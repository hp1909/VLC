// Copyright (C) 2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
// ALTERA_TIMESTAMP:Tue Oct 25 01:47:29 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
eds+Sr3YRBkwnPaHoZeU/VS+jDgeHAQFSKBfX/+rRqlulYyVWQXOlRyGsd4UUuga
wgb4f5rG8vGjWsxspGWXOSDLWUGr13XCpKdPE3mST+TdO8qpvzRowc+fz0N01Pcz
5T2i5ASm+0+qxZd9VAWu4MG72F/lGL2UPvJIl3zyK5Q=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5728)
MWUNCtRH8Hrd8qhtGJgJspZf43uK1+1c3aiVvllV6qI1BTAblPhPdJuw0kMgD2L3
bcef6mNwjx2TZQOdpaK5D4lW8Hj6MBBGf/M3sKNP0KMOVr4F+EILzzIQnSKdr9vN
mxhjVU0gtei3BVUZ4LO1AcwfvN/OrrT30MCdDlkSu+u2Q9BtJhenm67l6BVyOfC2
8g2rPmmBPScEy9leIJ1z/pxyHK6vzfQoqmnkljnjTjBHfqd9QJobLudym2I4RHaf
SxQG0xAUzctWqjTDSIWWDaP7gg3GOMSuviFlkhRJ1Iz7tP47xPFoIPQYeJ433qDj
J8+eUjiyJnx8VAgeApitVh/bPMNB+qJC70H+sSw7a3egC24SxJpNaHMcWhOtAPB9
JElMnFIbdmpygumMuNfdh2EiwNhZfkHDSOraGExosb6o6ZNjK6uqYhXAxHzqBIjQ
SsP4dYJTe5DI57BjKlKdWR2Hq/8PhoqNodX9UcmvRefu4NEYoocTlXqlP2c5CQb7
I1R/lyFiJhTP2cAnyIh6lcGwG24mJkQwbj4OwxtIkidOiQpOHYNJPHoOeVFerff+
ncIg9M/qJp4ABq6QCQ1StKHr6padbJYLaySNfKXLDjadrPCJg0c2gJ4jLJ9L4+QI
SY42ZmjnCshrpaowW32Tdr9REvbiIfokxjcfeFk58iNZiMX9Yvb2EX0n5Q7nOv0d
SgW1TRc8TOUuz0mkKOmTnF79wZkHuiSp+hLTk9mGYA+42RtvsfnRWS/8C+K7DqGn
WfV23jHiUph+fFwazNLs6cL2crV9uO1Xs9NQ3qiqRJlT21UBl0e76+0mE7Seu6mY
8KDwhZLVYmJsnSQjsX8MqgjzdobEfauwD5SFe88Pz9i0dL9ys2g19p/xVjvN2F8M
SIJoYiUxTQFU0Ewmps2ES57aN/NrucseJGIGyMh+SaRlxovD5JZhvWFH6zEf8fkH
aYmgZY/96O3/+kAn1C4B89lLXjtiFi5BQDB0kCnDHKhWH7604xTN38OZmQTfhwnC
J+YRHtBsFO7NuLcZeEkugjLQTuTPOiGaeAnd/g/alecYsudRKnJtcdjMwyfKJVEb
H/yV5hIUK9UBUaeOeksWfgfHkBieys0Jsj9NAf7Fr8HztCcYSvwb7iwVnl8bHCLM
FSGj/nF2LqY3k5QcVUYys9iXYq1P5PKGDWT/8dSFH63IqZ4VZZaJZkrXZFt/rngt
93X6TW0J1+CyiqxKAxtZp8qG1tqwpGS+suGGa25aSvYUJQfSWZsU9oLh8Uf4mYRp
ZvK9qFHN6qd8i8iQK40OMJVfze1dSkrQOvYweDAGxu8wUfRE3nwgNkN0Q46M7kut
O+4fJMBuM4vFYECMLT/FkGo/gp5FYEPq7ESmyTKgtlpuGi5Fc0BeY65G4jwIbZn9
vKcPETo08Cw5p7aSZDFefjrtaSW7QD3XAA8MvAZb9nsbQ8N3Bv9OanhVeXvs4Gky
Uo7Xh+ZGZ4NnH8YyIYd6h5eISSPcat0MvXrt6im7j6Lojeqla3qSeFWenndUs15O
tkwsU0FNkAxwD6CdVMMdqtkorTudpbTy4QvKk/Va3Qzl+/3t6zYMoZ7Fr+scAXnu
f8Y78mjGMgCJYNBoF5fEWs1TVrcAeBsQczGlX4nImAB41scBIVXdRAes4SeYnJml
atsr9k0oUbsTw01UbvK8sRgzsDNQ95hi1s9WzGI0MrdBXHAm8bC4AKKCtYfYBaxh
3UYKM8UqHI6YyVBBbzY5ymOwJCQ+x6vkrQtD3wE8fi+Y1QjesKYrwVceNiGmcQNB
kzOzVgKm0FJt7igd0nE3MxvvM22d016zZyI167c4OFkcHDwZQnPo9aCRn/VhWY27
6cS0RZ5fwLReF2lH6eute7QXbMYRXaEgnjpSIXJT/HTUWoEMt+X/W+BApUcjM2xp
p37itpyIyaRMtgaHVdSiKpJ3/fI4l/ZZIQ+AmuWOGHeXzeAVAvUQeKRVXuQmIxFm
1bL46jRWoimpGabm3jZlSGAR9mJKNKdEYVjdcFEylho3H/ox+Tj0W9Yf65EWCnYF
kJXTMcsdiLOtXpPnBVt/a2hydVjhN1uNebC+UApGW3F9UDRFmE/DnGmh+ZHYxJHi
6qz7r4hAkJnoaO7i/HIT50g1Kxi6f0xEc6hjYxbcUAxMpNqcu1XuD2HO53qjmAHD
HitjBS6I/1KqTzAko6lQPNn/PFjUCIROaUzyqBpNzu/RzmEuAi12NXMDP3b8xNSM
hEsJVzQbOBi1m0D0239uv++7pA8ZXl7O5qCj3NNNbj7r6ForLSZZcFamhzTdTqvV
0Ybs5daFtJqWX58CG5K4AJQ5KpwILR3q+abkJzQVJ05SZPkeossBkQtRRgcjhvRQ
+NPueX3VNEESNukU8l7Yjun4qQr3pVQw8zADrn3DjXA5a6lCOU1QfgrTFDXFxoiJ
KGMnu7116yNTKuQrfw1LLhEqSw12n52nYVGoftCV2HsieGi1FVukRs7OMJA9S7WJ
t2mlx4PBzeJm1Kob8y4iQCnClsOKuU/7P+W5y5C28ReYmv+XGytVU7NF5MCYinUh
tft7MCdpTl7PLqUJtmAmGmRvJCU7/dJJgTkP7SHhqMOA5C0xbOnN6zjzTp4AHOGt
BLHmb0BaQORmVM59Zaa3uB9/SEhh7gMXysMdlMBRXpYgpRUD5gCDn9Q9nd54LknD
IV4phY1Mu/mmVjOiISZTq2HCmkOd6kqZPQ2ZBqulPPytv4KZVrIt8nyw6xXBTyeh
be8kqOwYJ4Uihf+j7jIjNhC/p9rS8JVfb2WUVCH6Ux8kQ8odC4b8evzfFuhaFDV7
nMcUZpXpli9VJ6lXB1Vhb4bxCVGTIkt3dNiaoyxlTTvuA0kubHCnTepMz9rK+QS8
rJDzYAI4oVwWOu3AW4uA4SCBNcGl0a2dc7Aykbwr/WbIUPUNe0LhSqvbw94pSbUK
pUgHknxJqvd5ou8lsoSXmOfzoQKzvQP2rK45Q3H9TOypWEHOFAN1JD5NT9XRtW6U
sPMceQAISTSRrES7rPq5dqUHy7dMqqnQrsoWw1+erHZzhV4KXBSeb01tOU7/gNMB
D3KEnZN9nASqdm8hjFRgCtUafBbLEHjDqUH4qEHk75tvkxlLRfEk0lW9l2GWxpV2
i123Nl5/YMvagfMn+dzzHqnhquSQsNjmVi76/aLlIe9b1HjG4Q1EphNC0fgA6n68
8SqpVcKGu5Oih4+mYh03QSmh9umBB39ddrWwSPIfVO357jsABIxD8e3d8S5OX/cJ
qt4r3Gd+aA0Yx1Heg55RAa7EfICJsXAFUlyIBS3sipWiBNRArgorHHKscpsceVua
7IZCE9tAIOvOD7cBtT7HG55J/fTDZMmtnMBtfKHMZHo0qAO07WVwqsSemr5ojcGQ
o1gXeKftSDUsakOQGHy4CnATsJGqPGXx7YF9yh/MppWIMFV0NfLzJ0NwfG1BUdMc
RGerxKKN4Zl8xAuwbwPpYv4wRzgviJSYhYyAV9A5Qq9tqL4tYQ/uS+tVuIVy87Cv
54AEO+pYr4ULm7YQ1Zi46HLkkAcFR13v+OaJlDxSyUOc+237gk0vgYusm9XoaxVI
W7eaeGLNERoKj0a0c+vr3Ous6JQI24Id/C+TIFfBeDCCgNSJchj58EOd3yown7dp
wUcF56b+VvSV2DLgpV2O9olz/0GgISRLuE2wPC73JKALIBYXoAvfOgCpAHUW8dtL
3Q2WL+3tgv2/r01AVyuX7KpvrLqrtheNPM6gMR2RqeKa0fFeyeopoRlBqEELw3CD
ZM0NrMBQ1lOcds+Xdm+asnGq/R8KRw+8FiGvsIAuQWZecCCjQ//5vdJ/EeFz4h7e
/Ln8Iwu+cXPLBavWlG36g+86YJAkg3rFua+fpkyLw/P9ZtsI5vLcazgXq4P6ZN7r
xSVHGfT2FDt9G3JigwscbHo94dIXlRTC4g61+wq8rK4YyEw6FLjQfZ0TpNL8Fyy8
E24C0XSm3A+rgddPdBoV/ahh1nZvI+e8yK+zgbPTxX5F9IWYdONXX35NmKUKzVE2
2uCsFiYLnFTBRlBG6SB8JKAkucbUoOshPKj+3bjJj0Iz7h1PFg57QBnek7LBF/V7
g97FsWjHSM7CkDZWisfH8B2Cpu2aVdgnW9wBaV0Qv/YhrjzMaAVA85TOGw5deLBt
ZUkULqLrTNLYt9ljPe0oTUQNC/YbNpbii0jirQiNGIqt6lz5EvL6Ggtlmm7MxzeY
Nx0Iah/G/E49IbdOsPy/ucZ3K6kJwi6T1ajmG91l7hWDWiQr8X10nennDOY+Q2Me
1mUM9ck4OLwmTKajyDdRvjDNfmVqwhZcahOz1VyahJxWUdRHUdu0AfYlocSFJKUn
kqUoxYUeOtx5/OESOc/T/v2IgEN8u8PcrkFxlRN782Ij68Bwznoo3uM/pY9aaa/Z
RWEMe/3I3Sw2MAxs5TqUGq7rRUAVfhc11Z6/8AdQEWIBsP2TnUhtBVBcnDawKeBH
FDhUBLVyiA2ENfPfyDrJo8akdhwkX9ufeCZ5/chJ1yGCurgRLoD8i/5fmzUrWNoX
T2NcrLw2Z0erHXoqi7dOY9+i2k0mqUTlIz04bzxFuCSJvFyeBzK8B/WrOiS09ZVC
/yfaqlFAr1N8unQ6gDMz8tOpE2t6d2LPaXAz+G+rlr3kd3N+hLTDh8EdS3Wxz8W9
33ee458uw/Px/m6kzZEXmP5uNB72UdcDcPure2gp+gKRQgWd2fMIRRsweRv7xl0U
tGPQE+36Yj2yBDQQ2pVsj0RloyE3C2SJ5Sf/XSH8+mBW/3Z3eKAdvrheOr5Ssuzy
dKrsTU21AwWuJIFnESoQbCKCQHSUL1trFDvsnM9wfzF5JT6CMWIaH2rmAGyiaJHw
aOABRtHRSX5czg3WtCBfmy/D+/wqICLPR52a7qqhoI8W24vD7/U3xBnOOZITD0aQ
FXRz559MfRlHXEM+fcF+sOVT44CEtY2GIaHWSA96rAOxMvcrxMfq6aUih1K7Vd+n
pQWEV4OKUi0hf1zSamRyX9zpwBmk3kynKzyP4o44kkU/bwjIehbP8mbYsksKSqa3
UKA4DvimyzY8yq+OBuQ8/5yU4bluNpcN8KLMmqAK74xj6kUcz90nyuViCVzdE+6V
V4yanP/MCcbX9hOUe3/3q1LUipeus2gTrcjkoag0KAWBvfVLb8DWu8LV4Zardzzp
0Jaxrkm4P8206klDIXp1vO3wREiIzLTf0yrDEUTb584duzqWlCI8h//RsoijD4Fb
bUVg1R240Wk4LoBC9RgRq2I8U4uJwTjEga7ve3gp+UQuZuDfiI4L0RVYy6+ZOMvP
iPMD/ORhc8ds3fSNHimmyd7LQngUCCSKiQl/kbj+LcFhp73+tCIEGDgIejxHCiMB
P/hkAbz5lxjHhaWgJqKXNFCX7OO8qw1RfmW24j5bsScfwNXiF6xT9xQdwn8sfQ+J
0R52Zlv9Di2O3trZgL1O0LH7L67kgx33LIappue7qLshZ9BwP707+dM1u57EgFkz
kbxEvsxP11JT0JMSSiMONQKGRNkIe6E1zLdyzqHymhadmhD/da5d0zTsOEb0ql+I
HEnQz1GALVnh30eSMjBZqWChaIZ0NNE6ap+rvju+n76RgZvHed8fH08ssuJNpizF
YePF1u/miwAc1nA2gPTc6iBOltPGwXYQkp7kZKCsa1ulNeG/+nvdndCiYOE3qPu3
5Zp/ieCKFobpIu6dgN1eHQpNmKJpuvQkb5VqheA/yrF54kCSltAEoxBuALn2UUBg
RUcvSf/d66rI9c/wglewwc8uMvt+4xtXXbgGa/c5RskFQkJ2bTvEUY3C2cP9mU+y
7/zQYazD2VYVLUnZPK8Vo2vTBtghnHzo4UZ19d4l4bAhc9zdu6Hg8uvC7yxDcesr
z8Z7P+h5qkn6ni72wjX6vdvOGzqZO8p4Qx0l/ePFPc40+mKEd0FY/438/r3TAJrx
g7CEzWutURtEzQAOLevzUrYePyktMbXTAdl9pcswjuudFdu6xF0IVp4hTlwTViaM
shArvGMwpt2Ijek2ZJGUp5jgPCsKwKZ6exC4+K3BBtVxEv9huF3x6zpivl1GpRHX
9btxpyYnh0q3akU0Vnl+MqfA5+VtqQJoz58qxRJ28RatfrafNr3KhWnFARnZ1Sco
j2k3X+NRPGaIyVGGXyM+GznIlJ/Y1LLMpW5kmQiwvNK5c7My8j8SEYsp1I+XKA9p
Ox0muRjQr1j85YpWb6LHwhIcD7WX77Mi1X56wHGGbv6nyvrcracFfIr3uHDWnksK
dyoD/pP3+2KzMJ+iShIlS1Hz09aSK/lx+8H7Ef8C/vgMkI9UJh5mwHB5b+/hzyyw
pXpEVtvNWakaj2y6XSdSQVUuXxBlVNwEzB5qX1yctvHxfzuW4Z1J9aZvXiXVstRP
oRMwwK0dlXFaDZO/usUzFr1QfV6vpa/wpWsTFMR32bTrNIco4IKv6xcdMRGnJmLL
80tKpeDiaLcsubLOWnqIFm9nwA3IHRTBA3e7OilDdMFN1M+NHh2VJKBBjfuTDeU3
y4mM0JoIyGQoupu4EvT1L8FDX900YQqkQ48f/128hY26xLLFEK/QFiySJuY23FyD
LY4MfrcGfUE+xkEGvbJ+/8fuhvie7W5VLJgWNBctbbzlLkXUPSrXA/onijbz3urF
miYPkbbYZc/MNk3+Xo1FsghVkGTiKu9M1Rmli6sOcMOEtjy4ZUcqnwQdtHRIklak
9HNZID9vbYQRgagRhhno/YkG0ig2s26vdIshWqJsBKZ2L0/Z8RZrrQzuHwRihveP
t+wi+aUEA4r5NCw6DzKx5mgxHi5AEhsu5bvuGt4pjD16nOtI5dIIDgJPI+bsg3pF
4zne7oAFAZ25CR12bmZXFenLfcTOvr7+zjaCplfw5PdDLHQUZGc3bVwgSoq5o67p
oPQ16U9v2wRUHkhEAVV0sAbe48m5H1YezpRkS2IgyJenX+SYqgmgs+bMNGZd3YS/
SrLwsL29NEFz0gVjMIg/fQryQ872LWdq1b+EeLdPdKiz0kxHN2TXVl9pUXxh5H5C
okC+MdT7n5W+3Ec98N0XmdhsChJSNApp/i7gqHwHLANk/UAYuBeIzzdFZURbXQyY
98DJwq9EdAnF84xdoCVO8WqRPl9+yVN2npR55GTjakj2uwqm1BR5HagoSodaWOGx
rZk9RvabfT2FiGhBaY4FxnTCrhk9GfbHGC1dKSSoOAn6kkG1ltF3kdpKQmLM+izm
sqWfArwGpUqPfJphKIxeat/qPYz9nfbE9zwuQ2sHa0TLyLyG83mNAbedxOIVqpKL
3rqGIEyd+/9btRj8bltypHkjqabtazLd/OKeMkQvfU+jc+DohchQxFPx5gNLn9DY
6YL5pUEKLdrkic0SJqZyH8oP6fmyPS+xV77eVi5672sN5pRWcfqfI8cptbAubV1A
G7LMFDqaZsJAxocwPXrEawA6PHEGZSl/BTJQlQg9g0qm9RMuS1WKKLOyCUU+XLNK
28YzJairC0jXyFvn/oPOyxR+w9I6OEJW9MhtCBGLvgYUftlJ4XnoU8tLc4TSq/Er
eRfk5sWM+EuTGPmUFCftkCJQ+LQtKuX03p/CXg/KRnkrt5vW2EiFDX9s22KQ6vS1
HcivJLZbiHJO187elw12mA==
`pragma protect end_protected

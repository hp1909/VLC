// Copyright (C) 2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
// ALTERA_TIMESTAMP:Tue Oct 25 01:47:30 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
FIo8Ybnxq/yyi4QvxB5F+SpZ3KA8V6xkToqoHyHg543u7nwr0+lbI0UuE4cmlQxc
mDAuXamddDF5G4GNrrYuyXL4YfMBf2lDE6dUxYcBfvdefKXy+R/HNkT8R0g25TRQ
mLIayURPTvU4EVAQ+dlUs+sB/nQr+mFR5o1dNoGFFmw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 33696)
vyG9CRtBgJPmY9wJgNt+CMhdrKVNHJA15q3HNZ/f5TkJvA3/z8RusWUDyeleBnFU
uASZxYaFxrsBnVgD4myZr00P1D/XeeZ/GAtFZ9NBmr2FcfCF5+hOUGv0Bi+a/poc
GOGSrKciBALgI7XcFb+OPws317cjyyS37Ry1632G8wCtqMnY7FYlPw5UbVlWXXCg
KBZouqPyfMb27yj//tdCRa4g1PY7in6Ha/xbOJvvrD00jzpf60/r18WPGqzDbSHQ
T3gyrJeISv+szU4C8NRZlXig4zEy4nTNWVtOSyK3FhklITDAJmj7jOk7M9iBlwh5
n8XgwLhVkzYxIgSnzuUa+7RU/Ep9HHz7lkHMrO3LZ1BqiEeNapXB3+HLknCxW9Ur
Qgr0DZKohSVCjU0M3S1RVOIhraU99Z8um/0lkXpTKShMPkUnRs/Pgrpgwm7ZT6R6
7sJnhXOGAq3lfQ0Gw95hIHdKQJ+riIYRBJ1kGAQvGC9oyvtd1U6krqPhNEqPTkU4
cXZhVZ3tKlXv+AmMNYM3y9jDINyVuAlvPdF5nK8OVPbDRbhF+VIG2Wqx5IyB6hlw
npcscp66iTMjOncfkIo1Egk7/1K2GLnHFFCxxEOOElMPi1yRLdTsa07PfGZ1ZrDl
YH9IOYxrhHkHsAd8VZPgf7LF3/SB6nUamYnADYObxeQ+UeBq1UTVnEaqZkgN8D4U
Ow2WGP3sTJjuHDBGVOMcvF93l42Z7E6+gnXRozoenHN6vnS2agsskOMv9zua6pbl
HimFnanmF76gKrYRqpFgXBHKk1WL0gj/YweOvniUrkiv2PzMeL6dPSQj3qYIjWoU
+3SdlJP+xwS3SjV/xqxg50pr+TDF90Uj3McyU0qMfh9m5PYvb0lwfLLLJ3yz+MAH
r4rBr5Ml7/vms0+jcW4iZKPjSCHhhgQCgKE/l8o19o3sPOSvEzcwQq1UlbZC2aLz
5zPaLilr9h4SbXbiIGD4BtVT2e51l25mxx0NwYxup/oTikwWeJ/KTPZYO1vKluVv
7MITDdQjKw11+3dseqEuRKyc4mavsksOJ7PeN3jEGPPwR+33Xx6o7De3vctiATN/
IIHY8Mq3qePU7x3jTsafeBivUs7IpSlPYrwcmyY+SJfU8LgGTeCdXwq8dnk+zYgw
gNGPoy6FIUXeOjuQdi/Mr0IS2S5rOfm+ssukCoAVt0I3fv24DiW/FdoCGsB5T7yZ
fx4E6BgGFmkOjZci+lvquz3F7V+CI07zlZZz3Dh5/5NfrtyYXGoGChR8Hyp0AZCX
1eHPXfcNs84usrHGonBvaVyX7/2XVHLbsL5kmzjE+dQxkJEZPXUT6bzfhWmV6xIR
ia4d1tgGmtb3acJQZpF3Sjj/WY91hcGHYn3ENVhriaknllJBCAztwxQ2EKS+hJsF
jua1AoK4OTrAhqJFF+DcyjiGQpoddfJmnV+5IVXnsjVB+EE49kV+BuM2Be7w+cPY
s+qQWM+K7rzf1OMPe76yN6gn3jfMZq4tgJlea+azNaV1gsmSCHik/3xAxBYv9dPn
ux/xVQHUy0I4gXZgZ+xkGl//nqxWbcAINRJ5OnZ+ZgoeoNIe8bZTkzzXaCh9TK9Q
it1KWWOOQtXzq19kwHQSqQ04rt9jm9vZD0TLqncN3mH3IHhYO8dLnSKLJj43TrBG
awBKOQO0ckOoCiyuEJhKZqU1uWPf7spq05aMmrqO84zkXysp79f176V+n439T6KE
cdtHnRe8nY9ccZ0idWDo3+5rbQFgDNg06O8YbJAdpwZ8XZNbYUhic9iTwJ6BeTxR
1wr9ZmMSpuxurA3XqRXP1FaU7SPzZafAvEbx9fjwZG5cyze3pdx1s43rG8Zvjzjz
J+SJm/MFeGAuCrqC48FzC/iUOgAxV9vVXNwX6a5o7XWPiY4gqAvnaBDV+CCRvTPd
PWwfvJ04lUe8D/cIQk9ju8OTrSp2VbAZveTa3G1EioZcUOKwgDw4aW8qWuTm7Dmm
ks2Ep4cPDbp8qwvxFwfcMtUqEyixB4qWK69aJ+CaoZoyuwOgs9XuGU9A1u5RJl9F
PXZp4CzXBCJYd8cDrTUzfwBPp9UTGfEwEzt7BPU/gEmIZ23qwBacP6eLERg8uWTY
0CEKyz/WKinK0caHS1ErjmydaGe09NpGWKh9V4nIX75odJRLYPqoKIy/IH8AMklK
nDVjGdwLXrNZs6Wigsldpb/csg1QvLY09638v72imHjJ8yYRqhGtZTHQpjuEaDpJ
Zlb+8Bnr6EElQjUHzCBHfoSAHCKZsCQaC8Ntzyw4GREYiNOdPv8TQjCHu+JVbFwQ
K8T8AfKCQum1TyO+v9GBEd2kYqJNbm0hldpcWVXbaKgKtBVmWI2ZY2MTa5/8XPPC
5jaZykrYkfGQ9F3IgBfvpWrlk7OpVwQ1Xn1MvJXRh0C7ji5n3KUo7Pn5r8hZb2rV
kH8S0YJDsr2EuTnfBkZesjcijdZ+SOHK3R+GgoPOWLsHSh5qJzDswkqi7F6fOYIV
/d8aSQvoUBF2ntQ32ZEWLibnWMAqQkP6X3VCSFgup0PRRv5SQ/CkfazD0sdqUOPO
ZEKct+AZU0AkOICKsEb9m3Xynd0P3LytYkyetaCScEfbxRbqtRNfdoxeW8oHyrwb
d7dGsprcHSOdoqgKWwy/d76RfnXbL/b2LHXbe94SqCW95eRDrpoAoY4VpbzNft2k
zoM3Rq3Fa9h7UMK8x8U7joIz57+uP5WsbKdjpJvf1u/zTIB7dSotTLc7yrTEufW5
7kKfBqV+xQ0V2dEgAZ61V1SlvTujp1kALSuzW7Qrj8xLDLQCSpo/wQoxBTP/iVwn
WT/KqPca9bwLA5Oq9s2nKdnLk9HVK+PZ2dk2nuQ4WTgJFr+h4hmtm2vaY9jbWVTq
aDzSqvjhmY3LGqwi9KaSYqTqSjj0zgccIL7mrOQPrS/MsYi09X1tqTXptOqOHlf5
7J9QNz+fj8B86a056NNgM+KohIRz/6Sur8sGkYDDMbHBW7cftmyVb804qEe+rlpA
oniqR6vjTnDT6L1adYEmsPjr+GWhyQr3xH6GK+6DNP+tRNy++CrPI9ZvKkckfOdF
iEB0Wd0aJzWHpzvWtMuFi/TBoOQ2GoOlJDYFMjIdXgeGVLS5PyhTwAZTUzg+t+Hm
w2KDR0ujIzSIGaf+4pGDlhUot7qk00MKQsKBvS4/Q9BFY82puhyiUhBMtPJsjmZt
T1wi+yvoHbfasaW2Cq95p7qHeILArjPgh+Eh6jXRNWW/T8ZjRjgEL8+mmOalpeh3
gOvxLb7mKGUgWHUJhDgI6vsVVtF+/VblfNtvdubF/NWaf4XfAK6grM7RsTfbhG8P
A2YiOLthiiyFfiGZOvDVaspUuFqrdfMMsNnIU9wM7iiaodPsgMKunFgJPftyJOTA
d+54vhp1/r0qoOF7v4M2VerDzIiBd4WYkiLaG+qTpLgN/eey577eMdcRzUJowC1o
MpKx6EogTnMIvrKp1/w7rMTjATKjURnbITPQJe8aBTeVKWvjBrT5vxItOLtbwbLn
d87EKFTsrT3Z+8KdfdocZM/oRmxJdFxxZUUWdi+OI56iJzXaBqHLjkS0qHqH5h0Z
dR+4pmVkdlm/K6czmu40ULAsK9+oGfK/WhuzGqq59gLV2J3cm2apRnIyCTSQTB8R
L6gTgEFWwbvzLu29xsYYPrRoOAuXj4BNL6SqTSUeJfid9zlki5ZaiRXYb3y9TivK
Y09+fcyizVPPHLlzCnfdjkduqVyLtfTvNkCV6FZLqRTrWArIK4Ty767Nwy9Q2Lmr
WuvF1chGhXxDdJO/1pV9ui7W8JBm+yrl25jYeDJ+q8GzBzMiCGfDLeUVUeXrhW33
g9ayWmUrf0/X+4qKbajXEdCBXircQFQD+xbQg6yyX/AoyAZT+t4iYkSdIINKFrj/
6gtsuZesvV/ODkHkxaQgKft/Clw9K2K65sqiEJBnwRKOwYYsn+S/F7EfEI1mYxn6
kOtu2aEZFu05Tl4xsqanq+i1ZTWJ7601hKYyMxTJ6fSuEesZMfm2chRUScEFqvSi
+G+aQdNxIVH0Smnp1xSR7HwIDZYZuom34dlhZ4o3tMWpewHikCpF8t5qypTSopmu
kZQgTVqL1XL4YBjeIYD+M8Ef2Yk72X2uYfDYsPuiLSARu1U+g/thyPAlHqbsVZzT
oSoV6Ve/HGLSB7o0hHI/UKielBvCFs32l8/yywtInHhmKLgP78J0zawb6Om1caFI
WZq9oKmVATDKDPZQZ8ipkImA7a0jymqzKO/VbrsnTC/yH9Q3JhdY/o781WQ1w7U9
IHrnT9B1xEGmrpHobx4vSaVviSbjpA2IZFCvSp+K1qMeSFZfpcGjuU4VTzoCUdqe
H6OQQwSF7r76dHpPUvjDd4rq/vTQ/YZFqrYP05rftUxoilKzboumCOzRzNRoR6vd
jEb2cFJJa14b7T6OxSbRo0HUb3UMm7Ipfr/ZbZRNhJJaErPUrGTeNC8l+5Zz8cW/
/u+nP3ALuyJZhi4I9h7QlT+QE6ucQirc+ZgRpYONQkYC3g1rX2RIHvvppDg399LF
ci4MAOBIvBZcoMGBi1NrkVsyqDyCgFWY6M9NuH05Fsw64t+d4kdtoRxy9kzFKb8F
EYHq87FwYsR+G8WiVg9o+DkWx1jqWzoJwMuXpnQOuSSVIQ97ymCYOgdeREqagDwG
hFUKZGdSfOyoz6I6xsy+y+3BEzaRWxMUo+rBL/0L4cD2dArNJhmP95a5E32GXv81
lLzzHXVc5YYrnrOYcn73iUCwKJ3ZSWokNTOPF7PP7dqD8QnAUv2F71GbpjcWwoYl
m33I5fDdSnIQxbpfNg2qai3L+vNhVOnC5rYUGb8DIXOnq9w/rU0VJEZvXBFZcp2q
+uyehGHVDS7aCyDjuCmLoduQ6GpfJXFP1j1Nh/kn7MEdpETAbsAGlw1z45E4Dj8D
+t1XCAN47k3KsVF1tI8RKxezBSON8qY+24NN1+gmSUP0QmNHdH076hF0iERk1wDi
x5S6zn/ZJiIu11X9fhbzNMfrFvK3r2NTGpc32MreXYY5OsiGhI+FvbG62rmlSqD7
DFiad6mInPD7O3dGkLGty0Kfvl6v87Fzv7unXT5eUUsY+y0GgySiAu+qJef93ID1
oPcBvO8wROdalx1mTVkLlDxBQIKn+lNYHMkrfmKYVD6t9to9fsAlT9mCOGqGMTPk
67eQ+fc1qNXJhIKTbQmH6gy4jgDXm0rh5nQySzoc+iwMGdblO49jUjL2ZusD+tQv
QEs7N67tijjaJgxRWABdVKCkaZ12qajAFFOHeGKakPPi+/ecoAK1FNgRw7oNQSp5
GubE0lEyCKbCrXl0cJK1A5+FKLJi009XLgUtQqAF2V8+bPm3/fkE69+FlVPeaVJZ
Su6C1HjnEiUTdp4NWQu0SvJ4zX9wMfFN2dDaP/6TzOSh79whWnrDJdD0tY7vtVw/
DNgA/SFzPdwS6JKH6lemZvGTWMlY1ayFT5yqTuTB9iojhLmJKU+/4ONNHNpo1MSd
KonK0zY4q+a5meic1+SEpDqwuL+wMjXVURQUP93ua0YsoxgleREn6cY65gu8kTuc
Vz1bDjvUdwwxuczxx0rUPlnbRGJYBnBC4MpSJlX2zDbHEpq+QHY+K24IEMPn4n1k
nnDayKRVVeAttV8yDDNIxC4zOVaCUHeezUx/xrPo4sqQIui/hnPbq3VBIpb2RLpj
Zsenc/gk4FBBIemIyhe/kt04XSG3DtToXaJI2Olfud8N21Nk1NyVOIyPMmYE8jey
dz40pqtVv16p831iSxGQiunzDQSmbjOeA2OE5Ex0qk8PUdHLrGbFHtNvidcsA7Zv
9ZGyxlJzr1EO3iwsrAFdzdEXSSOyjlOYPzZvpqKTRnsuGOvygtQg2BL7pwHzWA9f
2dgzAMwu2H9MmY/iM2eP5QJk7TC5Q4+B/IWDOMNz6wGrHR/4JxawGIBzn1+y9JEi
BvMfSDV9pWw1tpdmMN+Qw5CTe1Y4We8Zz7dD20rN1iaTnQrjpjnVddZxo0HiMTPK
ZjfOYPxeAAm+LCzFEq/xhxZtjt/00ReP27/gPgKscydoIIQ83HDo+6kg7r0VBacq
24jFEpK5OM097d3qCPCWynxE+9NtSWnIY1BEK2YQ56dL6QbLc+C3AGnKyKeom5Ao
S+jprzwQVBCbIlDuAubdw+Wi9LQqe37mWRJu7aoGe6+ptv3PZBicxWyHhII6Fl/X
pfLp5c+65um4yaqFqBP05EXbBhSYOYpcJ7RN17ZxJ7Ftpu66J9tN2JRpsQgqaDl4
Fvg0ahvU/rNbujyKz5nfjAmEr0aH5XN8me/MmKTvxiqWJK1eJFuKl/wL05VDNTm2
F37KIl/X7+MBrlCrxqyD+jrfTWMC2O0EK2LyYQlO79ClA/008bPAYpWHy5KzpfJ0
T1hhVis8utq/GkQMTJo9rvL+x8IANFkDjzOjYMrFbU4ljQRXi1GFmww6fWFmknn1
ut2piDnhAQ8yyIC3LTKiKY3ou7aFCIZCwxOQs3pDqpbme0PYhOQHuVOdJtqfNUqg
idywXTbh4zjGB95n7mlV3MtWL4WnTPJL+mh3JRr2y6BruRcOz/rdRVuIVOArXk/5
yvJNEfeAHwoXPisVXTB5HJxqF9NMAgS1JACwbC50XyPWWX6qmaLqcEJLuQV6O7Jk
MYZakpfPGDlqImQ7Z0Zm64xFclFrkUDXq+e7UDHK3sNyDg3/QvvduAntGdsltcoS
5Yots+8Bew1OJrhK4JePq0zoPexd5kEWcM3zEgtIJD1kieVmPNvx+qLBsIB7enKS
b6j3Q5g7vRXrjLiLLb37O3BRjyr1EjvwbRCc3/67GD1xZhnp153B5psx9fZ92xzS
tBgOnR8XEFuLcRqD7D5n7s+30mu8ZYo4u6yttGYW+rRRE+6APZ0Oa3fxjbDap6IR
PtGIhhfQTy3+F6HPwXp1kMSveXdXvjykZN8CCa+qL3iLj76FGYL2MnN9lVARtDi3
0WFGfqiBzOKfCfAL/1s4Oo+WDiEMzq0o25cAi0niHBKeuZslqi34N8iUV2UAOVOC
mA7SSq5+2z7KuQx522veLX4myDtwg+E+Ysog4AEa+1zRDQ4fh+QjeDZsH/ci5suv
cVNNnmggflVFTUzqKVjXkZ5Nr/KiiCF9nZ1YRJgI6VCsrhc73Y7OO4cnXnqt84gv
oozmMw5Okobs9e4eYoEOq9LLtJUrBYT3G1szIg7llBbKKkHI66aaiQH0E5dUWphj
i0ekH3LhcVsXDmQfqj+3XJBS1KVALcW4Q9FvZwbpSc1LR1pPsrjBH6bFDerm2Vq5
Y+lqG9TcPlniMkSJE7sOSUe3AI1kQLUT9ff7BiNuWPUyKDQ92D6/bCWsKIBsbQLw
t6tX+Hbv4A/IBDtcfGd9DhMh7uAStXlvF+4GjovObZ4bFu1V9P7LTLMOFLEna+wj
W6kY5NF6qjOBRt3HcUvoKYDqWj5YctV0fgyKQUE2jxIpFv6aLaYCTjVgQFaoi5tw
JYb1Xl40YE2m05RHhmM7sD92SQHlD+rOcouaR8N6TmEm19fKbWAjLNYWks1/rBfw
WVaeD5O5lS5JPTeW1w3yUs/XUzfacduBmUGuqMKBd8Qfv83rPv00DXOUxv3Pmzy0
ere/PX/8iWH7fuLN1475Dlh4IeZX1P24tWd16I5msRTt9mqBIKADjs0Mn+PWRzMx
5Kpc5QnI+L7sVmRdIoi2Ypn41xQ4qopRZ3URzgMx5KKB68JWCtf9wtOtK3+E1Vgs
HR6b9BqX0I27G6A17qgI3KBMFHdpO0dxZtMVxY1XujjcKyY8kOQz+wqbwuf7Us+W
c4ZNFtEodi9rOXyGrC/2HrMwjZwPsONFmnuKGoAz+VcrRmGadILhn+/5hW9Nhb+u
4zFAwitqQveesSdLxTSEka59hyzcWluBN23XL8hX9t52y7AC2hoXwz/2m+xx8/hQ
MYY6r8bhtkDRPmg39qP5HVpOmLkmc2T4C9rm9zuQIxA+61d6YmXaG9AIB/I/sjTh
xYtN5477uaOFPcv5sy4g0KPtfBEX/2PAmrWFjQscXQ0t8sLj6dy99bDKLSJuKsPH
hkPTj2X6bdJh2tlp+EgTLD571ZVItz42XMWJWpJIJJIwQrVPiCey5DimSzMhx48n
il+1JULRngXO9XuOhDX4ajMwb7HRYkFE8aMvnpLfTata+EUasj1TdLpjJ1XL+tP3
2LMinQss124imG8kvW6Q77qxYhWCpgJO9XmaPUsTeWJlOP9tb86q7mKvDwg3T4I2
2tL9UG2JJFGVxDBGenm07V7t90Jb+wBZo0boeYzaYr7E+SI69vc6jIWsrChLG3JC
SH6HL6HU63PQGiI96WLAAYaCEVkt8Je46U5C3TdbevPYUFVF0WtKfvWx7XU9r1Am
tIfd/I0YUcMtUbALJ4eBxqxt5E8gzEAjT213qGfVZ73FAPHD6g/GJrPfBE+aoL4R
JN6LDaACDEC2BR/uEkxsf70Zz0vUg6/Xze4bMAgh5+EWKh5tnuR9LJsrghCZHRz9
maxdZTIh0d4N1KA7cDOHKrjSRTvzZnyLcOo9jnEDxZm+XfaiTYYWqKdmiFF77lGC
H3+vzwsMKk6ACIv7LQV8gpukLMcjQoqgab9D37/a26df3BkVtogk8uIJ+7BN7Oul
UEnFP2JdeywLYiVzlMwn80QUcbK6hOnH7Wo5XmHafTiUj1qG2vdWU35k+wJVogFP
adSpnw1tAWiho6FcNDewnz2ijkMLBIe0aJEzhsQWZlsmG2yOHAEJtNevUjHEsh28
7s39OAWHznhZYzJcR3N1NLoSeWm/keMd2825ZElf1RRD/d4udQKrh0BPVPOKtJvg
OaqNHeRALZyv7bjSM+EBzFbM8mXOrOk9vw5yZ2D6yb4xjwP5yJqq/JqyzMX09PmD
fZOCadVK9IiucHvB47YFdYPl3DMwzd2KcW2OVXjsI/gGeLluLMpeC2ikRHfPkjf6
HWpzMwQTQIHmQG3HSO3LEQF8M6+4aaEM+1+jZDua7PVKsEg3dlmMq2Wk0MGaW54U
9zKC+ilMnvoKwFPSluZiJg2OGQZ7mwWGH7MGV8DH12CJlURJdWpddKwT1dljlTYx
PoNc7fWdeD6sVZC4m5ghJJPRGhwUiGy4EfLom5ct+LV8lX+OkabfC9S9JaRjZsBk
nxQeRyidc9F0XQaXq79VYTW7ptJ92hIwEnJGooFHH5cCDkGY5ooa2SIBDWx0gZo+
oLNBspbij/ttgFhYC+0XQPjqStUTPlDeLNcAYNLhH0iJwfYzCWtaUEReMU4kC0g7
raSPgbSqOrNCV9hdC/+H0GXjKKaknW/pef8H+ZaVcxekJzVT1qcFbOm/XJEg+XNL
TiMLEYxwE0x4x2LYJGbZf+3F4SFa2WgCnIzlOMULUbbZodF3oNA6wby54yeBe7pN
PYaC0Ldzv0BiOJV8lXRckarw4xfhDyYkphFRuPpY7qosLKnjDqTvECcEtRpB+4yl
woqR1tluVpThaSYvgvUNloiKyQY+15H9krQYwH8vWGhaP5Hoa0DnGZzRT5F+KI5K
ILDjQptO5OjTgdUKOZfBn9zH7ndE6r9PGgCPUPT1NWLAGBwLTnLsmtH7dDNz4UTA
Lx6EPcUyQtCCsxqtsEokEsRb5ADsUuWFsbg4DKTMep9WwJlCr14OBuMCutYnqHMM
nhhIJtrLZpVaQK0iiAci7xt0J7y9K+9EslcaB3MjyaYud1Q3hsVHNGBY3qie6mUp
ncvVc2k10Hr00fsKihCUrZr65qETOhAvQKIwRnNOl9D+fppJ4GgGzTEcyDMd9QEZ
/E499J2XfCxFskivtM7/HAJ58L53mKBnHA7G5NUxfmX3UDsXwMnhCU4LSD5DYkS+
WL0Rf156WtoTx1W/+/NqprC9Gc5213S2W39gkXk13OU3aJsaaqnwkEP1sv3ie3ic
InFfH5N9cAavdDFprIuwPdX5MZuOTaxZrYUvephoR6cHXZv+KjdlcaF+A7yH+pkx
tlXqRwe9L5VcDNeQjdaSWGrwEQYbcORvJSCo1rWorJ5V60BWeVE/kev/3lBP71bR
VcvMmw4gEuwteCthrV5tX6Ik+J9G6gB4HMjIbMfbe2kKaDS+IGj0vSkWoCaWw3Hg
pB3xX1v0au2tWdpYMGPJnlK2Kce8FH4DZmQj6SOPvOtCFGAPvkHsMEm4Y1RULedE
XQHFKNUk0L8FNFplwYhKQXfqACoxA7YLGFcvj7gjhzecGxinzoFZB02NnWhrb83A
IvK0KOOJ31bKbWIRz9DFlDSXbKeyI4CoaqR845r9Emjo9iqeS9ynvgbV6sS3Oqqy
wp19s8sj5gzqSSRG2yU/VyUKZYGr6i+ClE/VrrG4zyONDB4dxJ27YBbrVeCZ206d
gxy4M04Y+pZk0hWW5ujAmt+Z0wL4NCne5mywpFS8jAFzDWdhwixzydv9b3pOb5QZ
5gV1FNEzZNnaLGFHk0pto2PiwIpJnIg0h082c/zyWiFb9yo53uykGFsRwFo1qygI
+Mckjp1jk/2cDWxycdKhhIpQ+cN5WORxO2InucojNRxSKWS+/kfkE9qq2EFnRLOY
KMfIUYT/GHn20QkNeBLdy+lH0f09poqJjiuuNWYFiK3FyIrqOjUlIfiKiComEDSe
6uj0jSYr7pcHDOeUI4TvO1mPiMBnn1zR+v59t+2Pae65h+CNEdH31pOeNIDoearg
Bk0eZ/Pu5fL9tcYV3KbE5kuFdfRhVhbGDU3Z+VQdmv/ifIUQF6VrUjZrTwGg5qJy
WO1M21mKIHCpaFPkwg4kD1t5L5rYxxu61H37wsA0MD1Stn3G6nJRNQk5jmRsJHk0
3hpmaLSHmo9pxAj3yheckf0TfHcKtiMmFq4zR56uuZeoSzdBWUW8qAKBjbFgguM1
s/SvmCfxr05AwPw8Y5shkI//avYje+0nEXr/tQm8ZE41awlqOFUEgw4/D+Jmiw8J
/NNcT/5hKqfARebIPL+MI6cjIZ4UTJLyCPSbT4ftoJl7jel1hX8bxe1Yc07tcXon
L5U7EkXcONZ3kWQc93TJzxcr33/155R1fJoJKRBy3jR+KOrjxAR+nnxs3Q9xeAYV
kwSqJM3gOH32sCpjDS2jLpQkqpBkacEHQnd6rkmkJRZA3amSSgmOkqAUCu658c32
JNvwviyQX1KaHRvBQTB5AVbmKpVh80AovlZFz2kn8O2DdPZPIRD0FN5Ut2xMSfjQ
N/czdvEb5YqjhymjQBg64WX5KuQiRPLGeUUDlmcDkBidJAR7AcYfMBzhNyv7ALwk
ok09X/AfGnYKJZOJ5iQioQ1K+omQof1PutXaDG57CvVhqNJOL1UAHP0h19GcMlGt
JdUiZxmgdE9LYpZ19CEpPf1Q6/wkjZkTJ3b8tFHcuTWpa56pEjQ+eTtsCB9iiVDK
yDlZ+SqqQ3oV1n2X7dRtoSVIbEyV11EYmniQbUmNjUiD17gZAvOSI0ZZu/Aamxyq
Y84QofJcj6qKas9giDTepp9+e90iP4esrrOTaOAqDKLwDsnhEAeRf+3F1d6J+4Be
j5NFXBu13OKpczwyHYadEZo6mF+1KF/9vL3x4qy7xs2Narf6JREtT6szT37EQTlV
kUA0Pow/Hv9R67Oqa+NP3cG+p+1XzTiQ762zvWRMwwZvVII7Guewa4bvF7c2yNcB
1p+s10YL8PxCfYO1eLR7oga7NEr41ejxR2oY8LZ5C8kyiceSV98lBUN4NrTYfyAB
Sd9E360IB+bORea/38h1xUYmjRVwmuw3vXsI2qWvHyMbCuKGWEFckAdBBtdkF3gi
iotRuvVM40faHFiGZtHpxhVg2xoIU/p9kdVXG6OwdC3nZpwlZPX0Xq0CDwjscyes
kUnne1HwYxzhzSgKpfwhDBJKFsQ1R1pwJjO5i2l3+73YLgFE8ihtFvo3ndAr5jmQ
F34uMEgpi05tp6o5I4oMfrCjQw+QBB8Msu101OSqAp4a9xQ2Y24IsR01zhmKftCD
BpAzjGG+V2u2+OzTpdn/W3p8H8oS4Vl6aF+ZT169vdTCLpWVKvd9mM1yIwqcOTnO
1tX4t4bphHxWHY5DuDjNnpgwORP/fX+wl8lv+WYEvQRoWBHXy1j9hDeDLpvQJJZr
Ud75lCv/20cFDpMpyTTLVUuGEjmWL4OT2Wn7auHm7VT8iKD2B17MYdKTeUOy72n3
Tj7U8sauakOvhrR486+FlINYxFeBxO7ZUWuSj8lQf5gfRZA/2VPES3BoPBvmT/qR
LAgmCYpbo8rhg1VZIwe847IHJWUwWgKVSnTRg5kGvXxcXx1Hk48b0qIHOFZDX+ZY
zDcrZuODlq5+meD7kZG5yDWIGa2TzW+dZeVbTCdAPFNSylw1hdDdMt99oOY/oWtf
KyX2wXZNT0OsjhqzPBJt0zfU9UMlP9wNQ26Hpn+KJeCYtqth0GyPpgEHrJ/SxqZX
CEbtBJU816lhqdkd+TmBOYo4G3aVziI8U5UNKbFe5yz/vojRbBY0Idn1YQ3WWqNV
SAOOOUQij3zVvmMuYuWHlo3+gtmgfIR8VY828zuVJJRar4AMKyGT1sOz+/5v7mzN
ZHQ3fK2Yq7rYw/PX2u1URlyZ8JjNTBmDEErlTzBFHJ2RFFcmP8Rr6PcJvgBzmhjG
tDB4rtZPg6QyxUKG0fBhv0SMLsaVZUWePi9kH14ax3yn6lhrnoE6LCx6EMrGk4Mb
9Rk4ZBiCHt7KX+Hy6RSQv0Co4ZCmOS41nOwphxbRPy6/8EromY+dWlLvaPlIZBYG
YBh5zkiozI0TRfqQ6Dc2qQtWEwIbHo+J6UJZKozPJX7IhwVtMv6aTVNhUMOduYBK
WamOtsFkzkRkzcj5D/1XJHsY8cwpyjZElm59Rd+fVooXRI9el3J8PXClHVct4wty
NQghJ4vQGmknQiVuVvN36O7lbbRtxOwzpI6GCH/vtpZeOawWt+G9SluwquWM0blk
G4Dgahb9joaF76/NGx5zK/cguXvW5bffa/gq1gppY3mgz4fxsZMLnxjtK80anWup
SrfZcfVodGMJ+lL4H8d78YRZ0NxTSZcq1j7CkEqZBfUhrOBcfJhow3E7zkBYj8pr
VdqgEdKg+xbELLj0nuOw668AjAphytjNBunKNZJ4xfKdjOJL6d6qnfcAH/mNz7YE
n3QNamH6+E9Kj1FYZg7xUHxQsr7trT/ea2azeP4p6HRTKZnyOIbCdGrNUVp8wS+W
U1rooRR72twvMDKgfhld27Xwo9T40/0Z0xXmfWzKS5GX/kEK9/Sj3wUDKnNdetkB
w6WvUELM9u4eoNUkjj6zGYYnwV5zopkGB4AbJ/YAvyM48fSbRIa217aNAhGDqUG1
6b1OO4UxX3p1aFIAOAot3Lkh/1iYvuWxDtNzm8IMs31qZ7rXmapS8mR+E2SJrsAb
rTWxnDe7hgZLUphpgZiq46vw8aCjQwO0un0t0ifPD6RHRQ98Ny5xD6MuwmXxJK7G
ccA5H/XE3JRExeViAJ7BlUA2/9LwKZFykMH5Y2vMzj/itpHifN0OPS0pTZh1ZvDv
wF/hYrzRLuRp+vnBZi2zBIezadiJuZv11zandN7eklmc149uqUY8rSg4zJ9+8SZP
NOtRlejVqcafMIwtgYiZjZiBvRI3hpi0WctkDGdJ4kD1p1dYHqly7BMEpDUq4hXQ
MFNoFguwtIBFNaHx9izSrmjL4QKDm3eYxgAYFo1fAihEnd4QxZkx9hq+fVj8FISV
0k0V3PJUlX2/cyhTf1ZAWtTFGVn75mTORwpYO4tQJlQpaQNJ210r52rETik9SRcP
GClhRVd0qej0d1wPJqFv4Mh237luG1FBuSeUkJdNRqUxeB1UOSkD/yu0kOOQeCuT
pxXFrwNaccBUz+jwqIlqpVpW4N9VGZEZmyb9WqkiyzcLZeu0j9kENUlM3EWeqfUe
aO2vyuBj3Ajz2QnmblLJxkHAURuv8IPYSRmKPXRPRoEGpXslkdGgE0AkLlqKv1jZ
vPVjqJFSe49gTB8rqEYCKk5SvCZxt6lG57DxpjONP5/ie7fkjF9/3JhOtIRr8iBe
pGqb4H+DjS1475t3NFMHirgsWE8nPJ6EZaVUNwwPxSbn+3urrJcEBkGBJsQGK4XF
9ApDcIIZJh2J2fRPMxLu0oJGP9h97I4KEoWFVIw490DUpL6kw9rYdYBPGWPQM3Vy
mY1+mW11mAj2lCodlAB0Lz9XyLPnmDouLXYYfE9v3Wy1X3sUCMLdZtmt6cgX6nlb
0jQUw/xo8JuoC+ohsQol2KCsLxVsNtFyPKGoUwpm8H0XfMTvEB41ymFNineu2SgX
P77g1CazMNkZ743dKn4+gSmZf/FLLY8b9fJaUJYGrsc7EJfZZFHPNm6wwz0MHEaf
/THSCS4ktfbg84rCJeVSgWnv5Qh9xRZ8C+BUUegYIep/NeREdW8XAue2DqEEIviH
+PCH5+TYtkfIMSPMfoC8NwiUcSz+MkIwocVSRaR3mN60r/qSW1GjRHhxPaqtDKAx
ttyo4npLQoVHaspoe17WkFIkCL5gh+uBg1GkP/Mko/T+ZZ3gX4SB6Ys2eId+RBWt
hi0MalwEMc2sXVKeAM+xwp8xFZb4ihHgmbmw0la4lZyOlpoLp7VMGxPGDf3OFND7
YBuYWTyWuhlkkeuesTCf2GsADSjzVC1WADUx1zvs+EfguNrosubT7rA7DNW4+AoS
K07lZ/GJLrDA3kBSB/kXEE1BZfxarjeQxKJ3Zni0A6w5VWP9NY0vMwY1bhj0amP2
iw6mJw4uJtWEtVd5m5ENxVqyUQ8Gs9l2KaVkNeWPOfUcKUAZ9cq9dXA/a7pdWbkt
geNQQiB9V7HPhBeOzlwBkNb8gb/En5i86mIRnIaP8UuBCkbckt5rtuJtcOnQ//9c
wO2sL/AffVhXLdZ4QwtYrSohsBxgOkHG+yya3BOmVYj/ZfEayPfDgfH63NOYbUOo
15EVbDLHi4dCagjbRw51j1djI/zq++Xo8P1naXqHjjMoDB/FFeOO6PWNYD/Z/EPX
1UBN9jTGojschsaKgzskZo6zk+dX6O1ahSzZRSjqr50Obc/eFM2U7PP2q4+LyLvh
EZNma7vcU0vlGMfvUIOk+xmAmhmrSwkVRqcZWzi0uFk+BVs2uk/FVJdJOXXK015u
WWkmephN4Dvztk1PWEI2lxV1ECNqmMOx5IWRzRRA1QE/umRT4dmm3B39LdNKlU32
7g+rbaTPqzAUGvgXPhvjptTofQ6aW3BBd/c7A//oJ3n+9+TGswiFwfaLWOjHaMX3
QuXCSCvsbILZCaSUgOj/rctWVz6yaZA3JIPlIREfVpzd481N39BIzI2idEJ2J/Bg
QjzkF9G9GQnyU29i5CE5ymyqXKKrIAlY/e09BwG0RNI7FxKDHjVnucnpyRuv5KYA
NKZ5TZm/KmkqQ9Z4vRsuB+RRpSAF3t995fb8sDwoTfiYS7Gl2A29xObwQuEB4lBZ
IsYUTtfokRQ+/xZDyj77/ujPM6Hprd+ecc9GtXKupI2Nin9kURPbMMYD/EcS5g5Y
7vBBH4zMizPUeT1CZvNrR59IrBRsDNSX68UCoqHkbYt5x0rSrjGjnye5K46FevmP
0OMbYPLEuKwmOgkv3t2v6VYAq9VgDTOtk5wN5/tnHEquOEsPzbcXxvK0f5saxOKx
+7iCsaL74Rx7KE2oFF+KBGSp1+z4SFBFz8YLguo9nAbN3Ehq5tutVgxSG3wmu1XH
yF2+kaj5AVQHNrYi9r54+bIK9ORg41DUb7ED+cqYLKAes5veicfhHDI/Liwa4PTF
fMG6262sq0kIIBF96Kmds+M6zQ584xHVL1GxpFiUHY0i/od2VjffIOhpgs63UwL4
56QYo9eprYWlR0wybwkG2Wbw3GCuHzY3cz4Go03lP/eh+DuNNodKLBl3PpOI0Gu0
67bnvSYiFauvd7Z3zoIHTj80RW0rQrSeAJ+72SbeyO2OZaEM+8oQynJ2+ZDnp0Iv
eonhaqZ+ZbbkdBmVn6pTXRHF3VYImNgBDVrDJl5hHm4sCOMCwYrGZrB9wQmWQirJ
1mio8VwmKC8UxD+9fN6FxreU9WX1HOnNUA8gSo9vLBSQOiqNnMm4odIxp7rUs/Q0
uQ9s/wySbTWgIqUncBj5bY2JfXkoo5TY8f2JfYMpoVYCGkbVZhvjQNZF4ZCYN4M1
9OcWLsS7chhVhMGosUOt8cgyeY5JxWcxgafvinWfVGbQjIELYohP/1AwK2nwuIao
bZxw8aaIr4GTYTElzUrxHZutmaDttWLb3mqBKPVpJw26GpScTyESMjlMvBpJfg5n
zAHBGaV6leh3gUmZJejlm91vo6DiStVAOOZWnkrNiFFRblwHKgrpbk3QWh2mG7EA
FUa2SwgQRMbGb6rYH0Jc3IpQDCEDDQQZW0Jqx0nP3/uIV1VHcul6bJqrFMmWqdC5
YbnpcFSNPyvcC277zN5IE6mJ6UOZ6ihtmFPqxVBoJZYbAoNF2CAkGAa+7svMGIiT
i51AXxD1BotYJ9DaXBy1K1rQUgYX78Imy9c6Sp5bEeZh/uVDdwfY8WOWoJEsNa9C
VVNCW1wmhMVJj6dh2ZBct3tciCOGpOWM56g21KCZa5usV7R3BLy4fePTH/nYS6eP
3QP+P4Ms+szZ/0KfyiaSI15bJVUNuikqfBD0fabM5LgdyTcFBbEJXVFPH/oTJ5HQ
K2EzlRePxT8yg1vEqmY1z4MqLYzqZ5FDlAJHA3Ebozbiw22SD5qCULvxc+483+ad
pd+6Wojan1HtHYF7diwbTfxkZdySCEeMvx1DTdIQkTlS4r03Lm2ymKrUCe3CTB7V
hFGld+izN9uYUEXSUm+RU8cB4o1aW0Yv7wti3yqu8x09xIcJax9tkhVVg3XySvmg
jmqeY9auW/W1aGI3bFpYIt7PGxwoP30vDazJ7WhyJ2AZwVpBa0X1W2HDJcRAISkn
DLXAGlF2Ke6/x6pcbYDv+f6BDxtjX0746FDUEASBzwyqrm7nnM/wuYCSI6RNkJWl
d24PWiRW+0o3RXl2ML/ePPyIJDa7dkfjZ7xFZixEtgt0xhV3lcz0acEj+WxzhQcF
mRU9OawzQ3GPa4jQfAFbRA72SHTEtsg24MT0JF0roSxzs0FBfe7ODvckoK9fJxUF
DS2XrnabaWr9H8+du8+mhmHfcYsdJEEgtGJ4cnQxCfxkUh+aEF6Zsd4l5Oq6m0+Q
ZQ7XKWFGR3IosND4SiqQhln6rwc4e2Pnbu3usrwhCXtNGtwvM22Usuy5z2bJN0su
qH12Htt+k7RXMUqb5e6v1bkeFekxS1uFh4ko0pcFNdxdkfsPVBvH/GN7UZNPg4t8
vZ+fC6qoW1aScDBNQL9azeEsPpXiXECGa4KJoeez1k6KAL5bc9KwOU4mwb+Vsn81
8s+7buC740WtZ3jcp0CqM/+EAeQAlLgAOzwl8ZcMZSuGOv7tXzWsdzz9yYU9ZLUz
xjUOD+JAU9SNnTvPXBpAtGtT/yf7Hwvt4A4Qo2asiseNyYj9zyc2EwX1mqSeyznf
KSKhPFAFcaU8q3WwjtbRdcphrBFHih9maVSxm9cYyA/xUC5jAcqH/CWwd/9kcSTl
lbkXEADYoZ2YYcok518nQYXX5CAKu0pQS/jhAiqeLmFD3lRQpxRHK0NrHCm0gQX8
WYGhYJsvd8+KZ9QuIO75hBQaG1/po8Dgw3DCYoOvAo0KlKF2DFh+qZMNY6h8c89C
d9XvcMjWz8Hg7dunGs3YwWO8h7TzVFWrJvqlAHtWsf64fUc9EU8uo/nVPW5FMQhG
8ZCoHneCmjLzp4WMzS3qAqcHFmDBka/7WrRXKR1UsXOCNHx/CCePs4nVfEJIOM2P
sFcl4QB0IE3SDS3t4CI/hSXw85PuDw1cH29vuWU8g6Pt/wxcIBLO76OORHHgQwKY
lscwmTFSBzA25534LCnHlc06rXgQt0QnFDM8fRbKHri/dBVq0Wn5nb6FxgHTDzhs
frg4lAoGZnno3ll7A6Lm+roGAQKa9QKwCQLoLZRs1hFhpuQMAPbLY1rNKXNcDo7f
JeEaVIvYqjQV22R425Vh37clTbMuYd4T50MnwKFtRWMkdTwBU30PSK9DCDTMr1QG
jWgpSYYdx1QHUfP1ljSSvRI7UBlfsb/cpEUbG48bK55y/uN/MswVsOKI5YMl1jwa
WHK+GRuvAAYVjjCZk2J1sHO4nleyB0vgSCvleYsxDUiFdC2Vz+utcoZ7zTU3ovfI
9OdtOaqw3mFDSx40fmNbH4R4pGKmBusNcrIQscmQugpLJhXbtDQXed/7K99JC9RU
hNU4wkc7Vy2a+EQasc30lKungxp34ODRvPuah4OXObYNki9YpG/k6zEg7F2pxb4Z
ivL9hluUnsv/gFkqA4ndgEIDv4EQhyNPFCYRMVAPUhvpXt1bNMCKaz5H5312C13g
h3AbzGzk4Xj0xqmxucKsLVMBfwGg/sPglr9300COMEQt+lDcvOFtlPV9moOllP31
x1Cmv3quLy5cnFaab2cck0wpEZKNm5DC5qVmx67FvBl4gzfL9e6nc5qW6wwvRfj8
eX3NQz1eF9h5G3hxGmzReIam6c+WDp8vkjygn6fTMpaIQZahuV0zeSxuqj0ThWYt
hGZXYupqI6156ym/PsGAOG4FBhLpe/zs+iSG4YwbSZoqmSexrBNKQnyNkSmWbC9q
EPTc9lOd+x02NH18T7xePGf2AhVsvBm75uHz3lmqOoVfrSzSn0+8tKN1rXl6ViZ/
JU6zw3HbP3RCwkQcOW8xTyldxV5xbsu7jb5RgFWXgg4Kzvo49fgVNYAZ8hcjGocW
d0c9B6vNiMMshGpKt2LYdBqUhMHRnwBas0iPqMk8qQvRIylPmvvAfq510O6LU1EX
BdTkclnbkklkr6Wb3g+fG5j8UeRX5XXhCf4zgwp7wvmW+CmrTquXoM+EpFI7GPak
7WSZ0Fefb/OnubjHGJ/bPEPJKje4nJBU4akqW4N0CxVw3dkGfZSEvnzFdIirmx3j
KTLxiyWhVZHa91bMMRsLpUftdL0LfCBOcl0fe3xSLbiz0H3xORytLsjmlQupsVcy
Ny7VsvlqjnA2nmog0NjER10//SEMFM69SYB6wL8JkdVf/90K9BKv14t5qoL7Lywo
SlyKcM5SlZjGFMQBscCRXbaHqooqKIMPYbLjCkarH+vyTkENZJIGa0uETkew4WVX
r0Ju4gG2wSlyonoYcgkt8A1IPkObyHOW09ZLWUQNUIfz1XICRC2XjZDzFPcl1CgP
7tqChACXZOLAhBXQhNYyiwihHXbV7y5qZpZzx8aghaGzG3dSJkgOIYkcJq2bjGyv
zpJ34MtW+QSaoydKaAtj+/nqGhgDpSowGM2OwwkJ2Qt2o6l+vrfZ1/V4PGjNjCMK
W0Jfc7hARTxtZQ+pSfty9mQl0YCdrMt11i7M9Zf1mj1J3QvO87FJvDvVYEqU3xvv
NdLaCTYG4Dvay7ocsLN/RThnGjet3+mp0UVN6TVmCkZD/0gnqx9Ima3Ppz0vaDul
Iai+lS8lYgRCzRJT8hRll+kzH8mlFra0F7nJE33oyrktyuaptj6m04Sr/thgQRHM
vj5phQa8Oyall1bFRiGIusguCGlPpKOPw5I4wAjk56ErQYl/vrXuqyzMycCPoUr2
Ohyz0DqOzfLEZ+ypBPOVSe2K/wPwzWc8pt2TLz18zPmW0Am5LWjBE8tT8XS47oVP
Eg6nD2ffuQgQSlwoTTeQQow9YmlUJ1y7fmh2VeeM0bMQnbqo6Qf/1PD/qGY64SUQ
IM1qHmA8vA2f0/jtutWFnzFU4cxgrf9zklDfH3dHf40Lym/Qkideg0vmQ4TvNJ7r
/E4r3ozfvHPg/cnN6ax/kw4/oBrqqyDN6Cw8m3oW1gRy+R85kjybWO0Id7oxDCGR
giy9FWAXrB6SPnJ4n76rluzGVH5V7B+WNC+bjtnd5pIPFW2wL10YEDSW8+0MgTNY
1+jptaJs+nkIyME6fkEJNMVU1bfIBlKuV1zD28MB31anBBPS0EJ3ufGtKHP/S1ag
2r56p56ReZntVd/dzmhHha4XAl5W7+RzBmxGVsgWwkZ8Ri23O2x7Fb1Bxi+EeuU9
YB85vuUvmWCSSImPxxtjRGKr+t/0NXYG5sluuWhnsVwmFq3v72kX6xLbAXijJkv6
/ZZP8wNw59ZtJslNTXHlAcoQ5KvxAhngNQhX44lLt9QULXL0n5l9ctH28aUPIEPd
gFxh3yMlQbGYf9QksrQXdAg2bzQhN9N9k2XyouTuLiXWD9sGRqqaqhvXaLg9gKuQ
aQs4QdZIpkuOQQTBX4cHjvN4DxqsCtg8HajtRLxGB0BYwkAHo32kBtLNv6df96Bv
/J7dRqDw7E0LgcPTEvzbJttTQEL6tvOZgI/Jt6g4kjRX5RNy2fRHfnxrh65FWx2H
qyM1BzZQgGLYihHu1petOen4YTvXz241j507eFSYly5SCykLPw8dFjtLGQorMkMi
fHH0yJjqkc/jk8KBcHhGVAj0eUYIQJzzpeNVQV4ZJEfGqNhEFFWul39YLw0umJXq
ed6RbojuYCN0YuX4TafFR/UdoRX+ZukbX5/yRpsQkR+h/pTFiWpbdea1cKgoBwIb
fDvPPQL0NCfC0/erOWYlzDWPwuKPUFLbkztXLF0mgvu+dkMum//Kmf3z+SfU6Vpc
K8AfUalnFAfMa6Pu3a9KJalHcldMdSLyf+y+S3/gNDoQYiPgnn3nFR/PhvPfkLGD
9fb9HlgBWvdohi7cYuovZ6H3XzUt6t9GMQnG0NWjh5tRcjERIori+GiXCZJjcBuk
AJjW9L8map2pZ219SNAQe3U4hlUeiYVLRsu9u/dVCZj34O+PKTkTACazrOdG7t7c
5MPa//QhGzmcs/QH96JPs2fAcKUramkvgFjrO/FEXbnx8/NsWYdDMkmV5Dz8i4mA
B6HDFPMihakKUQdHzeTFzXZdAkwXkrto9k99iK3DW/GSgsjscYDWBFNstVsb3MJl
hpw4dmJSUodYCa0LiTDv9KP6qBpXWnK6Jpu/JE5MYiK+ZJzOTcV4L8ZNEkSeWwxG
tPGfJcCXhYywM8W+lnBWFsnkWJ26dMdoqyJkCHcRY4p4cTL5/CE8WAbI2Hr/nGB/
pIE/qWO1NKRJ6bySr9pWUHVrA3MKEMUS22YFALtG1Ql44voAOevjUptSM2hWCSPI
ze/9Ir6JblVwjnJrovHdeAFz01nWNkawWLgZFiuWFmTeuEIZBC2AWAdBMrR0Qoao
ClJGM7pZpBdOZL/OXocc6bcV5EI8Qfl3i137RREpI1n1iuREmce8Jwz9y447n83z
k2BoNg1LuQm0p7wXRmL4M1X7NLHKj9Vkfgry4WTc0hKbMlJK/tPq0ZG1KHE8GuQ+
1JfNbvXI/cz2S1UFQwsFasei9dLGd7bTbxUM0ZW8Yr0FJjw1VB6PETqLrEe5wVSG
V61jeRtbBaK3CNgz9NYqwXnqG6dKWqRIF1FuRQlr/QwGXNJdGnKzZN16pryKeHqy
8MZToI+/H00hETt3VeTB3lknpGENkswGT2uaBSD1I7hi2iu9xxTEiW4OW8D4JwBV
BXEBdSxkYuf6IFxbg59QloTJwJNW9zuvFIbmLy9o29DxjMiZFhOthyLpeKllffQA
4FrwONuNkNTuLSnFyl8EH5gJnjVDFOD0qFZ0u4urJBdfF06JvTxjd8/8GA3M0wNw
uMoYt5Uwx7GufJ+f0MZZaJC1CLXTm8AB89F3G/MDBKATnmjEwdqh/v57SpRYcJBo
ZkyYS9yGXVQ8+IqSlP2Zlt6TbPeQHSsecknDHmFr/jjcBwfvIl85F26/a4Yl1zNh
yS71NYpBvb3+aT2pZU6SO3Qz1x2UjtSwzywKwlUKW9obrXqniOc+uD93WUAZ+HNT
Z3czJpC65yjv4n26CdZKpLk6vx71goE/e1Fn1f+pemaLJKttD82Mvt2jmyfnPH+r
BikvjMtZRT4XLAoPJGXfmaMCPPSTpsN7ps2opODn7+7H0iUOL7uIKrnTEMwSidWm
Z0wGdDz9OKCfF06hKanBHw4F71QF/slSoxbM1mlnFfie1tZMDCZue4BFvSdPJEox
csh31tSb2dF9IdajOB1l5N2ZN8tHwfYWmWfhXAo0+e0t7A/1RBJg5ATa7RCJvycM
f9Ud9I6V7GTuce/9WigbSMeLjyxT3KLRri8a1e0sG4aMEOzp1Vd355zOZ4yJUdW3
26nS1M+pIThaxxcw6NG0h2mbWv+NaJtvRDC1gXWdQAXiqN/81Gyj+muRBl/d+sR5
9cTtselErZJMo3RgWArkXodd3NLI3VMcKB8mYGY2SaNmpUgdplT2nv0Scw18/ej4
3cn5jRUzBZ1L02awBdRKlcdyuMiyGCP4RHiURxfhEjmWnl0G2O7mGpZr+oVKtdcq
LhzTGx6xQ0cQvG69SxUNYoExyV1vALV63Tg67zEzjhqXi10JPonif4SvvvpwOIF0
cSLOw9tscrcwHrpiH87M2aBIRTu1B+hzOWVImyWfXD1IhrXfnTK97WaENdFyB4V4
WbyYwO9FtJ2TV+5E178c/4wkuzfy2Qp6A4lcNAlJY7aBqv0As4B0t/Fw1Wwxc/+p
olugcirq3tf1ccKHgAnib1g63P+4aCnot+96GbzfH0JxG/VxCJ9ngcrmxMUPyqJX
WYGrzHwB5qEjNBixvKiVZjLUAg+TRTkGWj/PrCMLohduaQjZX4PbLOTAEmN7GqrN
JYSQtH6qFxBZccaE72+aP5iYWYWdfyYsDvslntaJJP14r2zTIVQ+tCoavEVnqSFb
Ei9berlQ9PvI9WX/uNWJ3YAoWP8LsY2Tds7BR1fSwN9HNJ99a3tYmYxuKu2Qc5ea
kNC9miwGU71imVKa2hQWnfvN3Xbmq+HaVUGVBkCh8bDeKMzrnWG8tXc94uiCzSlu
wP7fTSIvQkR1I3nwTynXut91otnfBbb10mHEuBHmT5u5uBk52LzEGwBXnUXQDGjO
4NqqYW1/LK0nBayiznCDk8mf5Yb0QJrzLqGhIhmv7t6c6MVf77xplXml8G1yikic
Zb1b6j2btC+4kQCvuoYN6IcXBNLS4XnHAJ789/bAOV2tDn6e5f8yCaica6kkUfTW
EDqgScXW2LsWkaDdqlFe4mFf2T1kwt21k4TStggMUFPoGQJw+Xb//PIAskboEVSz
YrQZBIlRusPJa6V6iDr3psS+BNEifAa696WdlWZ0QbDKfsxtcuKcrj7DUEN/y1sO
jQR2S6jui+192m+R9AkSyo6vKZca5LKtmLBBDWfbI57c89BF+my448phxCmxqL3i
XaXIexo+SDZwMUig1/Z2IC9riEHF3Bl0GCBlS/gJP2JjDnwhvRfrMNNYm8eYOS2Y
/vPKG6v3oqKSFphsj9IzRITsogd3c29MsiSkduerUrMb5bYjapedbLxGGgJF+4d5
YvgqTrDHjCIuWGptHQvtfmAoFGdttRWupRjqTaeig0gavKyn1x2Gvno2tyrwy+60
N55vHdDwFCq6LH1K5Y9nP2Zxg10hCPcQox6dF2hKWNKTxQZKSEjMHn1wiHo15yJ9
A58MWONKhvyWa0aU3q5pffTcMNOCLDM8BZ+Bj917GeeXhLv6LjQmeU6YlLY2LQuY
wElsAebrS6lRI+Z5Rg8Qkaqe1zvA3qvYRUghki2hXB99dgMY9wLgi6ulp6XhWG3w
ZbBg5kL0k1zaBqK6Pca2Dzc7H9E9Hf7KVRCpjwy2jXsVtSKFxHuhm/iBEnsYNzFk
tn7RC8fjK9gMUFPNn4457P38DJyFcvNjPH7xt2FBD584t2nhlHiJsd9B6KLgdzEt
5Tfe79SCwBJ+AbdKUgjok+SKWkwuvFNmWE+QPHYXO4qmrhuzIJGTzPJWgoGlMN7d
9gZ/bd2yGNQ3766SKhaFS6p5Uc98s9D0YYPRBV2H+KgKgAxbgOZdJenkbBLcpCn0
CWNlr0mzidC3D2F1s8hLGALvdZKP/yhU7yMibHQqy7XQaTD7A8W10V2Zq4suMckE
FgNa/j3Q2t2j8TAqBBl9VIEYcLEZ6NPafRMggNymLw8CF3TEUlIw723LdnuEBd+w
RTLaVorNB6wwPdDzBi38obK2uUhW9g44YZr5yh6DWecmpjnHuP9TrqJGt0CleNRP
tAPpzBdGekWyyNTgFsGwLyGFCmfX/QBxMrEWF+TFHK8Q+Cv5vakirfCmkWuFAVGj
vLWVpamYUBo04ySHVebvL1qCg59tpz3I9wyXGGPtTBb4M//5O9zejQqWMZb8telG
sI3pj0ICTsZ2G0BO2RjCXG8c89xiaHUa0qFuEGl294Z85P5pgpXE1bsOvWy6ALuR
GP80d828KlMPS8zjDq3EjA4NkX49nzTMeBCV3YS7SZB9jB+X5U/1G5GgGPd935y3
mJO2f9UYhbq4b6AXjsCJKSL2g1mV19x3oMwRgVnVKkTbtwohsG6Tf8S01aD6kNAP
uL0weCHfNZkE1hwnR7LSNj7W9MHVKDBOSMY/45RmFVgiNEvIG4ICp2Tnrku28pJ9
iX7hgChX//Db2oeDAUij6l0IHKV5+jfngpqF4owYctd037PLaz7IIDTOGmFW96hP
RVt1We3ty5BIRd2kRNpPaoLXn2GVWDnsZJyXunO2WdOBkeTTl3N0tAi9hpwCWSbZ
eApXwIG0WinmT9AjDnfgpPeLanVB5Q+mV73yBKYOTfjfR+uxe/CKjJ2+a9xtC6gz
i6qqNrwK9J31l8OhV0wG6DCBGliuMxFNJiK/Cb7M5WuY+ezkxZDagJA0pAb/4qxA
5IvZ/r4oAd3nUSaYC4vrAjQiT8D9CC2SSZ6jkbtYlZaBc684ymDgnaCbscMVO9w2
ATHgF/A2h5hsF8FkfYGsZq1gl4d/Tl+C2pb7tO1UBj844kpaLXVzh25OUOq4DUn3
xYEj6Bg2W0PYcUAUoDrnvX0e9KyFvGUtmiPEmcZuClpgEe6geXtaiYywPnEBQWGA
4WrYJ1qtQqyW2YM+lpEGNiq6AC0MxLGKqxNx5/iBEsByHvSR7NMsgdRMp5BdOoV7
2Le7gK9YaIOAZaQ/JfUA2Eur1sjlY4Bm2Gpoh+8oUpC6m4H2g+6vuQDKWoMfChB1
bpovlFIrunwxxllm60aim7SDsFQiijf1FSYrIPPMovpm5QzKcJfb1LZ8oQFq/ANV
iUdwo6dOPzKCGtb/NeCWbwt8FcO3GNLkgPZeWMNTU3Ua8gJpLYYVn083D3Rxxgkn
PFbNzaVp4wAjhur5suzrAMpwEmuSC1A48I+OobcY8dvtAZp3Ayh/ELEZGyWptNyW
kZ7fl28dVXDdQkpFEPAcMekY69aUu+qz7HZilrlmy2z53bnUJtcd7jETfZtdJNmq
R+ABrkrU5OzeL4QvMEoZmM1v26TR7LqtGhqjM9cqEC+eEbLT8d7RnhPJFAog71Jf
xIAt0R92squ8iWk8SO8p0+3SxIa6bVLKnyHfSKxqRefvDMuPajs3xs+fKRDGglE3
kLFC9/yd0Ex+xJYUPjuWU5sVSMjhhordmCmSEPZLdMjaNzyhmY9sF5RIzXNiqjl1
S6QnPzdpp1w1v94eTCtQ+Y9cpQ051LRN0w+xQMQzEt5wSgP2dkZvCvOfMdN9ji71
4FDnzWdzy8ylKJM2an2knqAE14kkmnM0Lh0s0tshxBJt5enHj7MrFZ69BYmMRqDC
FbOPjVyc3RYn8IH/77gR5atSDkShNacY4JCeCMimk85OJjg0UP4xFSw5Qj7Ihu1z
k8e9zfwBZCzLC1+zynzdlcvrUSPfKPrhiDVGzBFHG1VS2Nf6yq5p0YTpSykLKfoV
LyP7IRcHV+YRKCFxYuUgMyOHVrEjq6wG9RDctqq+osfghGHlj05AX4UlMwaz1+vK
y0I3MsYaD3mHVjJbuVStTTWKRPRWUYmL58GqfBZMInPMIxx/X8G13gLySrD00wQt
BHLLORWQSeMEi8ZpAmBGOOW4/1wlF1o0fA6oTz8t8vunJEdxiQczixdcgnPOOB9c
OMNNTVM1Ptxau6ncXsNyP/1qkCRdTaqWhfmmF+e9/kLfyIQg3IphVbBg0r+pnqLh
gH4Y+TnK1ajDCapk8+htv2XFkuxD0+6zkmBJJtGTEuXYDvtlCVxBFc8UZtzAa7yx
w7CZO1gHh1dVF/Ijaqod5yauuzmKJV00JxmiC3Jz8yfHRat3j+khqHkxAaEwLDdn
HstznZjjw7A0lo0fLOEJoXGWLvIg9Ca7TVAGtbuowswvvqDFvN0+vS3Vv0hRKmBl
X3PFrNQYS+5jKN0wciEmu3TETQWeNdXEA4huWqVdwPvgH4lJVVAI25n5gdsnyVj1
y3oxadIw7+97GsTJww7QjolOfo4QgiAaErDHHXbtubsG0MJz/DjZw4crN/q7EW9b
zVh9VWSBfwCH1bA9U19QulfXFrinVlXe7zWFy80FK7NwcSQDpAiheVwm0yDIZtia
OsdFMzXX0G6pkddhdZVHFoqpPE35pjfgglideaWn+03HrCaDolnwmdROQFHtblmS
8YQc9H/bcaA0LPxg2W1OPb4iHL2BRNZLxVAt9n8n79ifX2rym9mtaQpzqmRxYJOU
IhUyYvdOW/vI6RJviXa5XcZI7wD8Njjj3mYoieo6ywNzl//J2Mt1SSWcJ6yNFT2j
AHytPhGyF+Tq1Ik4URw6xwsSJI27K0wzh0+cI34K2Tjg9iZLrQyB9a9J9Def6lNI
o9FtqhSJU59g+i/4jqvLaaJATToAXwBR3RumKzwR4IotYSjOz9KzVfPm25oaM6fj
Lh4Mz2FUFVPS8H1dVrHGtXp5MRyhXek667HAv1aXhFopLgw48XPk8iEM1v5/e3C+
foeqNtJGrsnXmGmZbVHFn8FNT8KMCy7AkOTBPS/ia1njJ2KpRKdKrcvamr4IjRW6
N8U4o4bM2x4RPAKxLJYor+XosPgiGlq5L1MQcYcE+pDhv1HecfUk64qD04wUqz5S
Erg2+1F7vQSpb5Rs2BlmFKDtLzdP/wvNWNybhadYkBoG0UWey+CMcL0nOryvgDds
62TyPsqMCcppK+RmtXV3lxBU5UaIJp6ZRNUkX1f5dGxulSoVMCez8cnlqKMuZUH8
NFNYewmnxO+uic+JX0RNUKf3QIlTSsH/jre1k/5Ql14nPOzp7ycT5TkcUzLz/O/l
a+fSQMONRNn2jN7Be7ZbwU2/DXvMJ/8d1soozbedHX7N3KnLx3dNzbPRpXdFsvoj
S7GGH40eWfrXzJMYDBFM8YGQvTMHRyeN9NfO0cdnkTpY/YjtjXJ6PO9eOf0PBv0T
fDEoUKrzMdx9JhinpPV1HNJU8EQsl1rHd25DJpdJ/OJ3NALjv92axpnphMTaEiLD
+9QXThrbXyUn/Tcs2+1zOXD11wa23AfM4rv3bJBvvnotkXKQWrEQBH7xdGtV6p2o
yUC1vfZAL1I0tcUZCrPKpyUr89xYdmBL9LRA+DKql+HL9pXplX1G5urd99A8ROEE
CMob56vHV+wQ0BO0oIf7QTfmA8Ge6DA9GycQiwPm2c9P0aBSJlw4yJ8BchCv4w01
29IdcWvrjpQCKEcqKYw+yBFhjVQ/Fi3w9KWccgjlhU5caWNRfZvV4yE2i2VPYR+c
pJDgqKH7uTovkDWCZBItx7zxX9ASVt5Ir3L/EDRSnN7514XSgu+AJ4nC7vbFWWAV
cJIHuBVlpFg096cMSfvkcd+p+/DhNr+kRM/Vj8vKZFFmCH5H1Sc93but9jt+0gSc
SbIVP+Cnsr6BRqfqnvC2PRYSiJyLS7V1xirDvCyUktpF//bmP59o8ZRNNROEztDr
VNsEWDxeEg6y9dkDN4rOwert4JoelnDCZvIse5dbezxofZfJ/fEBvw+PuwLQEfr4
OkvzROUWYXMiKSN4oWPlQlzNofSNmNxorZs4HpRo2fVTFurTqpmtsOSXcOplNoUP
s85tzDgH44xOnh4JCgXeCjU3W6ZbD1c8iy3O6bI5Dn3I6Y7i4X7DgiEj2Vv/80Ql
FrOP0mr14/gdgWz6dQ27wImvKgXXoKbLj5yBNnVD83xQhAKHNKQOAOYq/rD50rQ5
7riV5VCbQnEYj9jro/s6cTUivDNBUTQNibN9+d9qGuptewZNqC4S1cHeIFhPM3KN
OCDJqDwjKzHGRzDT53zXwhnnlHJKxmPiyxv0rTNem8N575wTxXviYtd+8S6khjUN
2uAzt16Tuo1rMmaklMHgxffmU4JaPgXnNOLYUbySokJOwOEjEjN5eA5rDQ15nRxJ
HHp4KJjUVbEY9Mm/K5QBd9Uj3/+n1ifNbBXOP/H1ORHbQNBL1mgQWP/+lFp2/qCM
ERaD9JjfMnKnWo0Zb4oCMT9LlCC2Ki61F3zmGkIy6abPx+oQYC7jSjr1wklBVOxj
YuKi8uuVpyixygQ82JDNuROLfin8bZ+i0su+qVj2yj99oUBlS0K6xYGdO3lHh9Ek
9UH8UI32xQHEpamBtQxxpIzr+0GEmkpq79LkKS8pNCY9hBeZ827cP2i4ij11Cl2O
sAQdWFGmdAHDID9m2PvBzjSXg+3mYtczeczCOYxDIGItYI2ZETUGdm9yv8RbiIDV
CA4jwFrgLWvbTLGcDUfm9Y8cJNCy9a9kUQh2dFu6aQoB1LMRrKQ1AaXquNuOOuY1
s0bo4hZkF+B+4gKICoGc2vb4mlhnK7ZrJ+xAi3Vw5WBbXiYu71IJx3LREkvWR+1i
lDJVAh7HsriGnmguqslBaMcl6xbV3H8fuALKVMx0ox/LoNB/aoHu65yxckFANqK9
od7cUcyML0hG+0/CqBbjBg3HtmYcRDFMcW+QqAGbnazIEd25dx+/Q4Yvk98wZqRw
WF4htBgmutVdrBY1ITKiyuY2OW2Sh4nuOL10F26IZMT3zZq0s7dZZpUWf2qrz30l
ZCW8FgnumXvJXNj26PqpEF/03bD5urRepvxiUbw+aM+qnH0DC6aB9ba0dL//ubzY
ro379KzSiRRGLYyTvvXLzOTnFyH2sidOaKZ6f+SREsFLNP9ptaN7OsoJ0/m9LZ4T
3KBsTzd0yl3t4jezbtGmGiQkjeBUtnqEXcqKHnx6URppE81qoFcvnlAjgT6BCIjK
lRxEbLyh0t6LNINbzbjwrRHIje+uiDSxe27lPpT3NVmWLvmVKCfURBx4CqYsaXaS
4SGnLuB1p6IXMOcx8/5A5bWVfLzIU7onb1LMSNxLQUAbWryqlZFT/ti90FAH1cpc
9M3ZrZxPHu6YO5gq9X1ni+RkdTyFnd8H6ERZX05Nf7d687jKKprALhiHzUH9WXs+
PzA5f5eTKmMbvJICQ9ySLjOJlpcbIzmt3cumxhm0QFdlkhK7yHg1civ3jOFoS3Xn
rWYscWyfZjrVmoQzXT1NSlVm9JPqP2xwPu6bGxb7sUwFGXIXtUBGrLhDtlRQ6lGP
F32w+H4XndP7K3RK+7K8564+z+77eS3hxzUEjNDh+0QG312rVCEQNweYBHi6XNlD
9uk8HjjjM74ONEGw7WQD4Y1r0kF1hLRaedNG3ybYPS+66FLduD/SoWOXGbKTaFLH
zpkLCP7OlMOwRiTKJxyffrcyUDwZ8OmU7x5QG+Ey5y4AyypANioPkvD4edhfDTcy
11/5BJQ7grATQ0RIqa/NNezm9tx583F+P6MiuBrzJnAgJmZA4nUSPlDZKLBYAhj7
ZKkzwwTdzm1/hLwRnE/JraQDa2ertAyGOISxVfmVB5o3zsqe0bybmGO1S//2jRj1
F3SvoPk1TXdDXlcmLAKWMWbT2ML2eBC91fwmQga5cFIGh4/5KWqmDVHkhVrt7SBc
raQBModhnK1DUYYB7NS84GJr0OxAZhtahpdZLxxoxbpUmN3wvLyzhKXgg5MjjDt3
GXwCwdRGUVB5OT1Iyn4KBGpo05zF/DQI+pZJ/6XhoN7SnbIeNGxiu9gA1OYj2/Gy
F1z2iXvwyZskEKblnaB3jCd3gazHB9fogQBN/7WtfT7X4DIQnYIDdFdTqmysRLeD
ZwN5kD7rxr4RocuscaVngTiJfrppda1tQ+p8vIDHnsxVQSGnP/uN5ANefIbIr6Dy
+ToWhxiG4bt6lbJrZOEEIX2so/KUEkWimF5stFYe/Fjm7KdfD3UGAYolQBxF+0Bl
EXJZbJlNek4wAca5BrAUs5+ZomVrZsBMmJLQsbE+IuHSnskgasFSGmVzEOHAY2r9
Ztn/t9vTyGu7sx8ez25ZcsVwN3vBBR7QnTiX4Y9LLMv+vrTxAn68uTV18pkKM7Z6
tSWunY16gGR/ZMSE5ZB0UNwclBvgYTmYV4yuRsl1pFkkZDNpByECc4wASe6Ymt0G
yswaYRzvlhYg89VQngCcd1TcOxnbKxJgrt//vNCmfLFVGuu8EW7T/Yagset5TfpN
vkXbwdVvUX+umHUES4FG9sbbMJSSLRfcA0UwgekpQZwOM79Os806/e57Mi4bHek4
/dOT8PYrcmdwopGYZj8ojGZz2GT4XU6mXjnOlmpBD8UJvEJgTjwrqd1YrD9p+Tno
TzFhLf3dYohIyTQgYvPoORsoTfxr3F0ZXbOwlB1Z1fV7xjOnRsAzXFDxgLRU7Qpy
3jQShjXnnXAAfQCuNZFyMnF4GqS719buPqxLMU/+Vgp9R7+JY6om/ZyAhVVoPBdE
IoatUEMAiqCF+TtPA4UFvbJUWDrmjhTqNzbtmhJj1kKfkIdtiYRjeUX7KEmcSanO
sccW8PuGty4pd0wEIkDoNKQpWoQljkF1tMVHHU7KZOV8Vc9W6ZnhztHpQmJ0TPLy
bi+1m3ms3OvcFZd0qcIbOf0I3hAjaxU6WMncnkuDcLIb9I4N2HfeUAzdzfF2MUTa
AHBOZP2RgdmAF7QXi/y4nRKKOiVcI0hRO/07Pr9KnVv/dvJj0nQRqwWrtlfIX8Ol
0zB6g5xLAwepBjXKDy/5Ra8S4fauePGpB+3DSRjnH7U3xwAudC22tuCuPhIrUBja
T8TThNn6TiZlJb8G6DZTqUHaQSE4H1EAc7onR91oyNxarMoNygpmMj82gwB4ptrM
NToU3GnuFjE89fsKl2xW3T5ZKksXZJpObv3nAq0PrjpGMHyexdlQzGWvBnNkfhOE
N+wr1lmLSY6FTaG+wKWHgdSFL5P2fxX5SWO9eOL/NYDmKL9op2xdiaUwTapeZ91+
uCm1+uNFLeDDkA7x2DzaT7nPJ7SyVqqsVZ1yeM8XaSbmF3Y5kSRtfMydAA9ED26e
PGVW/cVz9FbaWMJAYws0Gy7q6PvJhmYfrKrqAeNWw/eBRy1jxQEKYbEn9b1G4RCT
n/zPmN2ku05oh9XDXw9gi10PbdFCVheAL8B+y2ZrJpCtzxAoxPLw3/9egHYmFBGF
T9//f4HmARjl/ymkY5rB9F/zPv362WwfkneuMRaMdENAA4XrdesGWndasNiu0Y/9
RKTddCgJlzYr7Ud3d6Gyee/PK2Xlqb1pHCUpqa618HS6Iigt+7cEww6ezPu0QooI
0ks9d/Xz0EsypM9vyOWjaHGa/dOm6UfDaznzYXFIpj8PvGI5wmRxZy7HLAvdByfo
CJPyWdriB8uMXvYV8xJNYwknEBcA9qAg36WnUSQFSi0W+nIFDEeMsunAPwq5/wuQ
gKSarBn5YQXrGEgx/edr1r3qHeSfmUdWcwyAhc3gtPhPlmRrK8Z2TrJK6cUkmlX6
NbK/XWOqqpQpyqD/a9o8zNdo2IXwB0Gc9VObGUL9tKCM8rjesg914cS+i8Uol+Y0
OzjMOatImuBg7tWTsap29jxtHgPLcX8lKu0A6hcjAaIxjIaj8pxHJQiz5dS5/WBg
itxvgySp5XLyOxoNie/q8u5imsWCCMMViZkAdD6xR+H35wpQ6uTMxURjbHlTmkVW
Pn7NUnxbztv1/mPhaqoCxKYNHA7SXSw7ooqjMsNJbD/YK1H4zL8R7Sl78eBd4ckT
h/3DBKxjmOYp1xwT+6fBfG6t2pgDyU9FmF0XoG8wSzfZlfC40SkNmB/B6pQEe6VB
V4IjxCI2IBtFRZFX6YsqHqn+csXVHNQu5QrL4NzcY+A0tBBHeeUmnQ25LCYdI6oX
TyZdGs03nJ7xD3k3jQHqre9PeG17HL3mOfeCuH2b9oap4vo3Qzk8pdfGBGKWdg3/
mAlZgVknoj/ApRzhbocMcZriqjcqhfVfQ39yZVrzKf/uf6dF09pZyA2vQBy8cmnp
Ydjm4UfLa9EKTsTvCzvrUyYTgIlgl5WGPz5meyowZ/tpPdMfyJllxac1cHYoDXWQ
90mNd+ury6bJvFp7TSE6xQDK/c8lBVwbk1/NLEyLSdqmixXTYN72upKHERroAUIf
sxPF9ZdNaeubxqnhU9Fl9iZnqZrQ7jgmUmqVCFn32k2YLbMCkbV+C7e+MduVehtW
3d9dW2sDEoSDQafkO9wH7J2jK77TZ2AiFnqg2Ogod3goXzzf9yaDblMcbLcN7O/F
VHGcFP5Aj+dB0QoKsRHy6vqgvaHfLcP3zFEIXifhvLeKG2RGwaadGws3aA3HHeck
prhcH6cmw/Il+7u+PNsHHuSYLCemmrG1hr/xzuUxumOReEADkg8ADcZGHGc9nAHN
WGjRqgtxRIslFFtw+A45IIYiyia2t+xS4njeJ+OcigvMqBrMDhlv6rIhbzfWTv0X
/7M+ixv0+XMJQgxuLTrg8ovN8oRkgCGE8hanKpRafUl/P6GldzrkDPfKRuEMesr4
iTv58C5TCovrMrPU7SteWQ3wFtxPIc2iORG3NCQh5gR+QIOHfBBlvwYwfylPVYml
CcXEhl9lFOGER5iRKyPMYGprqwZP3H/WXw3A3PMpx9TomohAREjcCWqD2mJ+if7t
ao4FOVXnouNxbjcVyvZDPoVlP9HihKoX4KnaHexZ+sBtWuKBEibKS7SKbdHl0Ook
qqP4dPjRGa1CQp+L8grXVUVpHNrp8CR8hmF9tKMuHJ5JrED4XKPkxoinoix9Z7g7
hN1Rc1sYl3fJpnhA65aEzJuoyqnsXEC/69fNZQ6qacPl2CfqKQM1hxM+dZJBp+QG
wjhRn0HAzi2iYFQwvuYs9zAL7G8EkTsc23FnHXx5RF7/nD3IYlPWLMnFxeDm5UDL
3gtYCgklM1esVDA5LpraYPrAOhy/aG1qPOWr9P/nI1q1rYpI/tAnszwE/o8a69fB
qZTjFnFyasVDmScpHJPvcbZIkiw3NgwBjq1WdgCZwVLf1GpJcVluufOm2jfmFpsY
xclPXC/+8kzH3i9eGEGrhY5SlShdSoZCm6rpo+oCcd6IdUDE3VnaXWPp46lsPrVY
WpKnOYKpgWvIGzBv8nu1gqg1aikxuZxbsT53qtNnnUXJrZyGGqrQ80UVIjvXRVJa
U1KmNRExJZC3zWlYO9cVJM8yI9XrtLz+9l/8meggCry4lGg6ls/b8RmmxzSlHrHx
wq2Q6fSUYYDd+grYmhpRPACDkZk6d5T44cVyER3kmH3Zj2UBxLm83vSkvU+enFJC
Z3M/m8Uo2V6F7lWdTOZm6gmHVA0sBQNEPXttyth4xlTiDrFvZCfCVYW+/NtmY3S4
ibvZ0ao/PQe9qEIGhJ1dF00K3WhxuTv9a1wUQr1TUCrE0YBj6qvc9K5KhGse+i0W
TLEIqwmsdEU/d8dWtSAUZYoO33rFDaP5K/ill5Dp4x/4ZLGXsRxgIRrqwGM4y+IE
rYTqqOK4GBJNfE9EPxGuCLWw2kZe234PQfpy12TfoXH0mx61NpHozjZz8SN1QVwG
Q6bjR0rkUm/+dLWk8Fr8YpkvLUICuuW4XKsUwWs3jMT98Nr5xBVyN/dWLEXY1n0Y
CWstiel12w8UlIKOVAMlbbNbig4beQcmMZF/m0mjPcvgHL1hmdmEJhA+Cg7siya/
i/bNoVgWRNvkxRkeQqa0W6xoSHOwAyT5e7ds3TAA86XDBgrT958rQcEQWv2BQe0T
d+8BX61dwEeE2dPZP7NO4K979qBOCzvuKGaK9BlhQ7M5RxcCzhT4RjAEEqWRmxMg
/rjORC+/zDRwI8RdP3pxSPrF7ZlgWEpbmCPsXAhZOITFbz8GkD2qaAjTB2RgU9uI
JBaWEEMuKnR+UFH3B2SYy+PEpuLDY6esBmbUAUl6ag16/ZXgiL4S+9zfTQBuVwov
IJs1vqwAbeIWGQX2YC7x0ABnDTuZVca2LHRV7+EdpEMRA9wr/VcrEz95BZjo0Lrm
g+eE33M+DpQ+XgxSs8bhFupHCgIO1yvIwfp5yZdRGQ90Wf/COxa7zrdpyeHRjR3e
nb9ZTF45RA3Tzd2VysPJ27uQdIsVXRjTathfMgmoLB0NAGOc1Ht/nkiV+XcyN28J
KFqSsZO5lbZfABYTHA0nJFv3LwqK+VK6WedCuFZobay7yHH0My5ubyWLbHMzAXvG
voxMqzydJybCUOgsTjopsPnCI9292whlAdzuqU4swijCmvwPIThys9nCs1RdncGZ
NJHAlvRW0L0TE3c8CVhVues2txjGzTJ0dK1ibBkEy6RHrwVTOGRNObiPH8cjVLxQ
8lyUP7ehcbjTNkRMfdTC7CXLJoi2ucognImkj2G2c6PVwrLcZQVxP5rasDBHUm2e
WVq7ECpD4D2mSvBS+kcSQvpeWFw/eEDKh0cXV598I96g1TsxAuext2LP46TQ3qxS
55Wnggx4JeCn/KGD3SIDZafKchRUPdND2BH1+VRdPNoPmcfUeQeuf4b4izM106tS
Jxgl70zPKbeY5McU4E+lJl7i7PM5wwB2HviAIFvThhfppBo20d/96MOrKXkkgAfv
FfOTrCYEVAAwuPq5oYB6RzUbOYYQ6C6MEQmAU+rBAyhIE1hDtrBfdlnbjjAtsjSY
hyoad4I9dIXub1ji9OYwXaGZ1WWoc9jczVD/7pe03ArxPDjn9/J5xEe3nr7KJxs9
mIEkANHcNIvFKKTfQ7/HrxUw9zEXKYp+2dJia0GnBhGUpLqwaquK3VVewygQf9w5
N5HZBflIQCOD17Yv2CkCQdk/c2yL1Yy6OvvCrLOPlplgBgUInkbFGrb/9F2cBJOP
31eNWjHVWGuKw3J+0mMR8PiTbrrVlYducvIZzpUhMc1Ruwln3I8VfPR1rxAv2buP
cRjrXUmbyydpoDUzRWWwW0L6HL6JtbjS0/XQqItM+sc3Il3fT43bTYndVy10J/Oa
7+h9f3bLVF4mURwTV51QTug1YWEanmQQVwnLtjofLzRWgVQ1tbkjXe0b5+taSz2i
Sd89V5tkkESH3ZTErwfgEW2TqVLBfdGc7+C4xOytP9a4htC3zkEE3G+Bv6Kd6YSi
9GanoINVe3Geeof9PN4HyEEvy6llzaTRjck27Goy2x8Qwc8FcdMCBp1MzJcBZFP0
fIcgIYLrW2IqkUCR/NVAspLMnuSVhrYWwd7/rkPsrgv2i++78Krm1pYO9Gjq0Mwl
3dWASm0TCEDtDn0OQ4K20J1UuYt1F+wqsIS618lIVbmCVHUwBvuoOGdPz9yZtztj
4p14S6AzTUcTCuFvuqItVB99cx5kOEQ1wOO9UXV7iAIyHc9+sI1LIfoWGMu+4RYK
KNykSwiMmNICIJ8HmUT80ZwybRL7yDfnWb5rrVQ21qCxt6ilVg+zHxuiCgenRjYJ
3lTKsi2jBvhrBbnky2FmsQ2gDJQmpQMxW1ZzJ2Z0Lk8eo/Q5KSgb1Ti3bjDQkNs0
hd/XkfxkNm79IB81a159eAmIruBDadHjIuClkRR9laPql0cxftMT0cot9x+e8Kgd
cR/bN8K56bAcdjGqRkPpdDtv2Z6S3a3dsOhlOqhrQaH8ZTlMJlYNT36GbQ+SXr+x
liBADsolDwmXPMGBbB7YDxwPf/aUuwtQnrvdp9lcCWWYUgnXPcnrqbnX/KA1SQjS
A81HnMUrycjE72hHPGToe3hrj+dtviRcg9ZkdT8eEnFkY/DlrFT+HIjtXD0wuBOq
mISZThhQIUegZQ17ehK1p4RYKpdowvtjFH/dOrqAwYTVXRMVx7ACGAKQrP3r2DJD
NlqQUvk4/eJkZv/RxhLlt3eV6R/A3TSV3+qhgyonVoFEgXalnFR9bPhSafiJ3h/C
SVK7hl/koPUsqeXP1A161qGsUPKDvevrFxvXio6oaKz7aZXN9g/7C96HX523EM9X
baib8E8IHXmmkiDVmrfa3EWZ7F3TABWJ5Wf1IMJjAt/s3rPyXp53hQip6cZHNRNz
b00BeHjH0zTiT6moAcLMxfFQ3DxZpBE6CCwYTMdCyxEKGWv4JV4eNEqboM6rdNmR
AC8PHt95oC4QZvTTV8+hacU28ppcdlIOoIzdVQc7v0YWtYcJQqrafNJVWD8w4hZc
hEiACaJtsucZI6y9qydT06rBFWP+ZYBSrBlI30VhjR5nFJZdZvXdqitdTHE7FaM8
eWl8YCYgDjw9Rb8ufQd/o9lK96oIvjPGSPcLCS7JQONDsUQp6oOi+rsqe/j77LIV
RUtAsCZ3qNXc4ryznm0SXMVyHKPL8mN19LyTdImFTfVq+t3pCecYyy3cS4rl/Oim
KiIiYkRA7Us2ZgLW7t9PMKP0xrMUnqnDFTbtkYQFY7YbqOuglYr7kW6lGT0cEe/t
79AI/K3sTFqZ2y9I01QoYPwOHZMbK8k1vAxqWQVegAocLZ3Suxia40ZAo1+Aluq8
EVRmPutLvdE3xJhB3I6wsDNHpd1Rlfd3lF/oLTbK8mZOxd7AT+F0MbD3i+Zll+Tb
EPvehFcswNSJh0pdoZ3LtWzP1X/4APjfdwWCdBD+xK5aXhf3RPn6Jy3c9QkLmYhG
tNGrayfo+qhh18TtVVlZ3KR/YnKtbchJ0B7Y4Zt4WLXfXN8ob1FXn643QPCN8JiG
qqDgRHCIw5DBDDOKUF/UbOwyM+M70qsia7P0gJit3Je5TUo8rr02Z7xImeUA7RX/
rJo60k5M5ldg9LvXbi9blcZuw87g4CsHq9bh72kFn2nvs/iYErpd2wAXjWbJLJTm
KnI8ksqO1J82hnV1etwi98hFdQyxdU66pr3b6xRk6jZ5BTbc9fgXf3i7xJYMAXyS
JIezayaETJn3H2eaup3EPu1B6h75t0GEESayWZAwESCJuZHyoYc3dJX8MxOzdb/x
unDxRZtRUlDWgeMAIiHusfaIvaOFcyUBRGHuOHtuijeKjAiLLTOwiT/i+0k7yZw2
yX58Qt+0XQ7WUxxRIOvpF7qXHLmIgRcI3mAqwI/mbehdv07YpaeIP2CDo3xQycKZ
ow1xOug8klfcoxkUjFYt9NAoiQw6smgL9HfzsrFVr9Xso71XVhpx7T0TNjGFncNz
Vn2rDuUv4HHcnWY6Ccw1FZvgVLGeZIQSa8yxmePBCWMtwZTUIKrcvnHou4OpR1ik
5v54vJl2aQ7VFb22yjO23zswXB31obFR9oqhQDjNBYdQQWXg+IsMH5Uzy5YDEwR9
d6k7G0MWLrHJVJoq2LPkeW0SA9CCk1ZCHLck25+66EepGhYX5Op1UHXsjfogLNRm
WbS8JU4PRDvfQ9BdZK7J046XBYGpvvBBl6rJQhiwaLgjCELohbZGUDsyw19qvCOv
KPFQklNnidKmLW8zjHBhvp8pvCqkZq+c23IywGAMWDGGdpcibMSDD2plarvx0lhE
K63fAMHA0yhvU0tRauVSeJq8XrVbENU1gwLAZcprnZQDBptRpExOjL7g+uZBSvp+
0qmpRqMUhG20Yvreu46q4KbD+N0eOeT0ofT7Ok8q0zUAqy4MREwcvc0a6CAxH82u
bERnXL3kp4wom4XvSIRe05nZy4HUka8dydsm5JNnMecooZVoRnXSwOurQI6eh9np
pA6uAlw7P8V+q9FlQo2QWw/jAALaJA9BXLProC4k1nS31FMxxozJLBksn9o0y9ye
fT1FP2rtOhTYy1k7VfTAKPqBardUr1Sn0cPVjgTyMqceI1JrG/LKw67TH8WDumDV
aPWoMPwYXeUes8RjETmlbf9BmpfzvG6VnqxIB5kaDTDdeuG6F4FeQiCISxwny65F
yMUG00+kmVGVWnqkIi6nmoY/HCI5Q0NMQF3wMrGCm4D5qSrvBTsmSaWQpBwQknem
5xVHq3ZMo2ozeFLRp5/c03dN8tEVOqDib7oV8epFUzvFfgQjeSJWuWqbNTBTwfr+
85q1+Bz4U39Qd6U0UnkCdhkQATdAUjNH8DMashNxXzl0f4ZLdPfFmyIrpGukdd0i
xhC8XmESP0tx/CECwkERQ4iqHBag61Ptbah4CybbZatb+fEy5B6bMnY8jeAdbLCB
qHw5y4AfiLBjLVqfL2LG22qBntI/jIrkOdGUD5on2M3NGOJytL8x0r614oNkZnpn
Qq2p8Qimo0N3HP6dPujkHUuHoHcVkWQRshQI+RNVRZOivzJNYZf3Jz158naIaOhC
UK+o7P0B1S3dbh/VizALuz4OxXWNhSZh7bQi3P5/Fd+CGnhP0vYuPlEcq0XzCcV/
4hApSirtV5/fF75+EnBhHpSDByHCm/SMhmUN+Ty50cYECVppQq94u7Am5SDUl7la
OZbceHhL+O41Bj5twkt7bERbZiU3whNdJrqtzRxAFlbiz3ETmMQ31m1PyV0cOKAb
YjZk6aYr5mNA4WNrAEXOQJosNgrw9MVfZOxyq3b4i7ZF6j5vAfUTKZ5ZMmKIItL3
Q/hv97OHwb/QxbfdjwG9Y+2DsPzhg978qvpWIp/BBRHNu60J1OG9Y3hBz8uTluui
P3eTIGtIUnWwqL5BYG/tzVtW98noXzvUXf7Sl0o0wIVwHdzmlvFcWAd/u2hB4CkM
02bW+APyjbM18PpqXl3MKBi433iI+VaH5RQ7ilNAs5UYB4ViHvB8TATqTfOcn+8I
jFKoQ+xvvcfu548UGDAdsWzd9HqjnNvwGATljqVex8EvCW6kuI2dIMMA6e9oZ061
mbsaV93x98d1lSomrhzHAHiReTH5Z5TQY7IZ7lFFx147AG5AbDq23fgZSmqr6hu7
pHhY3UFzVn/SquyKLBhn4T1BHNS0KRHrAuc97WYX4LlrzlX/Ug2uuuJAGaG2ve3J
usiJqpIe3gy8tBq98bY6AOjHSNZcsLjDYGEVMKTTezMMyrDYDSkob2JPcrai15Mk
SqiNSpnPZhLVH8nrZxiUabeRTtKzSmACRBsKCOwMy1cjaVAeA6M24xE2b6PB4ltp
SC5ZPHglHFndKEw2N25gMuilTWZ2xNncKuFpd1PvT3vA3AcX0KYWNBP8R+ZZq0IZ
51zMKOb1ii6MBSQX7JbKtvd+Zz96tedyPk2Cs8Wsk9ToMxmrOLRYGPpHw1pBGbU4
+0y8HzO39/nFMKAyLLfQKOYhzPiJRXhseRMxh9jFqd/FvdiW/KBIRAhXs02RG0qC
qEdolBHXsC+QftEEI1eYX/PN1gQq9+Y0epm8OXB7kC3MmhnXzmrMsA3ohTPLFyIh
rVq9GrLV11VeN7SW9v6o9+Bg4nCeJ6lfuBPNOZ50bTsPO2ntPyOmpJJ6lMP1DbPO
7m33egL06aU5/ZPlN4ueS4/J8xEyARVArwrdOewTiknzAuBnMD1fvOsofL+72BnU
C6nrXKJSaO2u7HkHN+blXdzI2BaIijAm2L/mLoIHRvOiZGoKRqRM/4gZdIyUi6TV
FElNhweefLID6wL92YpFMPn1S3R2P4xux3vVn6U3GZ9TvACKZq6Pufm7x38PeZ/B
0y7D5hOtem5GV4QscAnFOR5tfitVgqtPXIopKOGJCb94WPBnevlozxbaZVHPexFs
3p4XbUTyeDWsQQfUt0/OYlqmF4hTe56Xwk6iITeHIFZM/aGDm8Cl2dH/1mB50Kcy
QUhnoaQKZDmIgrqyL4wiY4PUEv+ZNWlsEyVkBIw3vsHN1BLq0Y7SV40iFMyK5leD
j+u5aHdnrNl86E89aX17kjmN4Ot10YTeFY7PvAmZo9uhzzlWCwbrN59Ry6o4FpPy
i+KH289MT9G3xT863MKZNo13VlvteNnW5gjWvNOrya8XFauMIviL8R67jgIJ3Fht
dda/QKfHMZSRTqGLGQ7SBusICB3f49WD4IU1svbBuc4Fk3XyPSGdI2m+Z9vTb7ef
E8uIIjF3V+aoFp6yynw5tHXud7tOxpTiV+wFELEQUmSOgtzj9ugTi9Wczn048LF/
KPXWSjS1w0yS1H6VHbice0ei4kwJJaf9XVX9GRAukeo3L/bJLg3zb8OqYzZABD65
ehSHSuK2nhKXZuNEzEiuzDH1KLVW3JtrzUfJ/rVkJQCCFj3KckyzmLJF9qRi/93F
N5GdvObP1EskffgZC5BjAeFBbZ7g3o7YWI8zlasNPRAkMsnkQROGt0BX+SyqDoZs
ezMql5YGqa5hrllzC8VkdvIPDUBLHrRIDgGLr5oKa/0j2N2wtgfIBavqUQvKtA5H
h0cGxOSfipaR9LvjBBNlOxUFjQVQdkU52NzJGXus1SjVvNmJe7rOubZ/eIQxmOvU
/d7FCOt91l6C5KZtiz4Mn6rEMJ7BDYDCDPRmmyKwt/s9+H1rSPFSOcAwLSpJVez0
xq9sp+dFYqm6//rYqchk7fW3EkeNkxxY/gHH+zhl65FBlxypW4CY0ixnykwxAK1c
k77EFYeDb4p4LG8pypIPdni9iQ2e0P2UJ+ILcUTzsd0cDBajs4CT78eHQ8VuGofE
o29LtZDW2mccKZhBZQy5607YbIwb5Eo5zMeo8pHlISiAbv3q3NqjjUJs9y2Ip6cl
MfcZRy9Zm6/MKZL1EXG3Lyk9vazRRCIIQTnuLdZCPqlsKSU9O89TXyBcQro0u3Qq
tmFS50fy0AhaznNbRuVJcHjBUHmI5sLIqVnsnLlSJmHhAl9TzA492JCUcQsFTLLg
ZtQQruJ2oC4Q+ISXCOXb/ZtEfRIro2Op4t6gZJcA5LmRtklplkpMiaeGZbYGFI4r
+OlDjSGNlfkutkwq2paKcMUo3Q0y59u5pVEbGxHoyHRy9JF2NZeHG5eagxxOvm6N
mHKnUTNZdJXADabTl5sevhYLA/F+Ssghj69lK1MQqzxhxgjmMYxEp4WN0FRotPGm
2pcpFfi6y93YsZ+ZKsXvAVZzdPUDBTJZy0/o8f0KU6UVzV2pqXAdAE58G+lP4v49
a1ZN1+MCB7nEoxJv/pDllONKSG487DhLvD1PomWuwOz7ReO+rv86wx1Y16KD78Yy
Pz7ltaQl83dP6Wal9H4Eae9HSORkxfz+DLs3gisfXE01+poP8JFLpyys1d1K5NfQ
2scEIQbrwBza3ANhzVE3IP+eqtz9OGGYxnncuYOrLPJ48Wx4ixjY1OC02yymWCiu
PWDF7rQHVMEf0YRzeQAovGFkVjCrZccK1d/Nr7BKOtzjnG2A2WeGl0+2iP+6gbK9
luC36QIHsa+/90h+fLaMF0+Vg8kqMX8M+tnU5+0VBLZCIEBFE5B4dOM7TS8YbQhg
SVsaVrLxcIlx6+pGP0AXCiELQIi+q6rCMbZrVke3alDixCsPXTUmMECo+ihASGSP
W9yooDIOt2drzZ1sYbXBNhB3Eik63Lr5udYnjlqAGWK6ERHSfX44kdAb+6z4ZDuU
8bKh3fGvOKU07kQ9iqcg0l3Z3LElG2lpZu+CkJhJq5szECsupSlbawKwpXXCmvRV
90j7L0cdAOhOIuPaB+NP3yEEpGN8U2jBsNZc7VdatudgvMCNLjl6iywafFANr/yB
3ip6Lg6b6TTY8EBqaa1Hp1bOJQrTXR1b/Lm/uIl6W6esQvAVq7uOoAlDd6DDqtgx
sDnxSgCXeTdnALtGIZeiak6X42pkMLmhjMkYeVDU1BRBanIqBM9QdO1KvywXQrUj
WqHEx8A4V+nW52x36REmRXWBUiTj8VfICG4pqoMd9/BG3bNsnWrzzw/ucssEn04O
oYKfnKhudMpLHa3L/49hjlbO7FYzBWH9i4Hi9JS6mNcG3HvU9jY3FBdn3tub4n65
n1MpnG8fUsF0Sz58CnqgzQZ/ICDJJMUwoTRUjFlRwReS/y4Hz1M584p6z7OCut0F
SziPJscTswhin19IX3/noXvSV9TXwZVr6IiSrHu1IziRhUWwYxMru9n56UMNv+az
dXJCO23gArOvmXch+q3SEuMAQAEhe+6Pk7FU0zR/7senz89QjBtPZNAqLa/mX3aU
IGi2QYeYSyzCK6lcB59wgq4HT1pA8jIzQdIw6JGN0FSlV4j/mWuDfUk3B/GI7l0W
JEd1vb8xE1n4chig4d6c1119aTHTSsz32Xa2wCXzpwQMvyX2w5Sd4XX/WKPN7ehY
JS0HKwiigLmkWGuTJRLHY0w+OxUArv7JZ3ayFDro+2ku8IZGzfwAWmi1e1QckwQu
n1S7OjpA8V7/klzVdfCJdDiVHlEFoLlOpN2WpeY+x3Mm8BHNj1jMlSabz3SnxGl7
ACvHE0T4IGgujQRISSwZT/4D/f7jpYWfAQdESAvsCf9CQEe/Aku59B9xSyrIlDQP
C2VM6tcnW3lRP5S3d/H4QOxBSsuTTuiOPewPixoUuYbIa2pq3wLsgQjdYSYKhEre
PAfR4w6sjTaR/qTVJjTA5GodkL4BGOv5PoSYNB/R0AYHj3rbk5RAsWxBU6o2qdCp
/LUkdn2dyLxhS/95StuQmfvuFqkCu3yeBVSIKd5aMdZLtqd7KM9fx5nRp7vbFkDV
jJ3dtzk+tfgGc+lRx0haeLffgjZzSu6Q9xqCE4Ewd5TCPOZqQqzXj2b/1x4llRbn
9rfQdmNUO9s+8J0wXHhzsBxw2l6iKcExHWwe4IXy1+1ecKjAlCPg8fD2Ke5mSW3n
n/RWmYhAMC863aRqYP7W2gzolJjrfL9zbuOqEYbMT+NskdAJXdUGpqHzLRenPfLC
VaXkGFr8KCm4vwaHUr0zuCrHiCzV0/1sobGXS+Mk95GiM2zN3T8vokRtCLBDeM4s
AVi4p6eFi05Qk6a5hwL6QW3Cn6IOYC/AfgKm1o7bT5rb/uFzjwEmdLcSV7hPfxqe
S/18yL9+I9iiyJqwC90Ju0iXke7Tno5pWsW7HT75Ab0pVJ4gmedIqlIyg8CC8oLs
BEzfCLkgo+nfntlev6KY96jPLJ7PQZTPNzXHa3tTJOKYLKxEme8gANYjqb1m2rdo
zcp3bam2m/BmvO/9OhXC66YPWdGqofN3PlLyMtLPJ8FNzq+KLk7Tqa+pfH5L9mig
inWIy0PTCAHc+QC0b2X2Iye08Kmca5VmlFztHocESw+WJuQFr+NNDjB3SbXWNR1f
ZWNPe9qbiZ952AlUaYyHBV47AOZhWJruCcqBOa1JCBGGpawy/zjT/4HAxAINMbEe
u8YnUG3XObBNe+4asm3jVqF+vE3wb5RsDAJwNGRM8DVD1jqwng+gPSxlNN7Nt9xT
M0/CuJrw+hoF0o6vJSGXypXUA7yEejAN01FsL45PUdjXeIC8US9QNdzE44iozJ3m
M6QkqC2ontfrADLXt8PMukDietkz18YHAiyfUi2zrZ6/+tpsWGNHANl5fVFZDxmQ
jd1H50KvfGvybvxHiRYeUfRApZUq6YWepk+3Y0TwoiIaaU31qosAZxAYPDB+EtLf
RDwoPPy2iLw6Y+TkH6Or8B8NaxdJB57Nc1/1XzvEA4SfeuRqxBdvd8aXXTQYBbkd
WY8Ihq/DOyMF5joti5iCtYXY+BjomgjLpcQytT6na2aO2HkfWIAZAniJsAVEkR3K
8VOuzI03v0sY0222jh6n3CgMH5rN0NzsgN2iz1MNs/qz0RdqxAY2Ml0NMYjE9xXU
w3vphC3msKKGrXOya0P1dD/yGDlD08LtVV/Urw/EsKKbjMeeldl1HJATBvhkT31X
3i0+m1IcISE4Ls0ieiZSMdF3oSfYqd8wdk+UCQ0hgBiUKQ7ZH+7/yBQv3iZc3NH1
j9PhEX3IUfV4CRHs9EP99JACvZtqXPa5nK/ZUkg5FqlwTp8afxuD5zJXLrUvwG3s
rFdhKpYtzguu1EBj7aCZZBduGFgWEMNj7I1xqArFLr+svKpZPLYCckZcehkZPOi0
A0aVI/a2OG9vVmbBmXs1t2ad8QjuBukV6VBa/Xr9JmNKnUus3+ev/XcgBb/9Zv0s
mI/mmjEu8Nn+5hlrJ1hm0FQH8AmePmzRz/oRxmK3pv/wWHbv9qKGqidmgiKllEHj
QwTH4/LMk0I2F328s7U18aNNb4CeI8CqJUhAHcENqH3XM4VZ56zjAaKT6lIkHT0x
3GAz8tG0bfKNGMBmdcwuCMFO5oXhYfrj7CeOpM2F+rB/Dxs+aCFcAwl1cQ0SXyj2
GS7QRcJ0e672JFbmFPXymCqAt2n06QsAZhipThUFxVA0c2dDc0sBVLu0VomVzFIT
ow3/+9ynbw6HMQmc+OwpwGrnAhCMWbmCF1y0DXp+FE8CHQwvYuPvqS2NrX1lM46W
Dpavoh3vWu8C9HRXwSIdDpX1MA8+hY8SIEy46WOiRvBjLRQOkYrHcuzBpoBpEzX2
hyQ/ucgVKa/5DV2mveslV+pSuxU62OlRe2zuv7kaeIfenzoXhZ4KR5trM+c5TGoo
IxDf4vEGq0/0+iQzRnGBbtNXuV08yx+pXmnXRKHOczthSwq19iKEQ+yRyYAJFjyn
87fAIcGzqWid3zFfbE+XU3IimiEYvXtBmuSh0UGsNd37rwgLK1DBxvQvkgyIIjED
WtSH14U6T5qfIKyOZ76mbmeSIdgFV4Or0jotb+EZ01Cm7nEkHH7nloGKXNsDexjl
q+tOjXRkc/zsyptxJqHBpTdcLKhIT1IcGdvL9IzTb2YNGWNsGObG6v2+ATroD2XQ
0ns6Xu1jHKe3armPx9TFa/AnM9fz+4HNBc17/CHKs6XHXxdsz8h7ptUeAiHh9hap
OoVnHP1cSMiolecP9lKGUyniRNIJzyeSGo5XpP2YPxc6ysOuxMS0bL1zLLZ7GZBP
rUL9fvDWTvUXe3cqwd0aA8s/jYYKf5QDNpS8TAHb4D8R9OomcPbMQC6W2xpz0cw7
mrQDJnDbDC6wnM/8+fYcBhZ57Wj9JQtNui92C6MNmYaxGwnNShFkhCA4irhreom8
w5Bhf3E9INcnISDxcCrsntembC8yj9/ZKtI9+oLx119Q5p5W9P96UTdXbjYwTdwu
/1ZrvwuhAPtFqYLEcsvZQ9URGLaJwJ2dxI1fwkKOZtzs+SxrDRBXwFLf1QXpLpEe
`pragma protect end_protected

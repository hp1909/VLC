// Copyright (C) 2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
// ALTERA_TIMESTAMP:Tue Oct 25 01:47:30 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
o6V/SqO4i/tM0JR2rCV6N/3mbX+/WS30Ntvy6C19YGoXOrY5UH4qCrmnI8MDFE3B
aaJ7S7mgxmy4pHjr/yzzBCNgeNqZqiswArpzyFTW3EQo0wsx+9NoP0dtWfYaOXNj
KXTnOwqnFkFzTU8Zk2HL0xZ+2Z/TZ6el6wqiyqzSqcQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12336)
RC7IuSZR7UqO5WxPepIq48qmkIr/fE3rLj8daoNUSXgPTFI22q3k27413m/0E8pZ
g/9VxETdocbY+/C7xYU61owYIoxSMAfEphOrS8VVE5xFhJNovQSMaJnjDiv4XFB4
ngccgkczVVrWx0SpfmQA2flsv7XtpD9BL7EXTuO371tlXUpk/UGZHGVcVcjxOAIK
+IbdYPEDTaGRi1VNRwz55PK8ZnYmgilGvMHIvvkNU1KaVF4mMtlnrfqnJxl56DkM
pN8YvGUy55mdpD563wYpn0WAXFlzfqlOlnqAtwREm4oLxftv0qUutqBNMceqhftn
A8fHRwDw9q9M7CxLhIFcgvO0ky8IcDn6IA7gaZPmFbmY5J65tP5NzI51tW+NFPUJ
wcyjLvbOhbDwX+TMibinpRMqdozft9NRQf31QmUjm5sjRJPATf2q3PkzciE/N6FY
UcpYWZxjpKEIPi0fnmuTSqtH+uGSOYANJBBa3/qRI5jnd84EzePHeUJq2VaVVLCi
L38mGJnZfw3UlToH+HJdaO7zEx2D6DnzI/O+XAzH8AMx9wuuyaViqcK6bmtfSHHH
wbcnjpRCCNTxTKnBxSlR2GqXYUCKItL4BOTBoGLJT6F6DS14MP9PLwHGhPoKE638
LAB+bRGq0nR1FH1WX0aj0BOq2lK5kXcjkBTFb7HxNVzhIrGSi3KuPpHmYGQfzWsw
7VBXBADI5fs2eGdoOE1dMOxQwwkG03L8FsEdr18Y6oBetcyJkxxjIvCqOSRGEwEQ
3mSmffH11NQqocqIqpBge5RSv0DkRf4qxV9/D7ra4Qx/v8Ix8ImyWf5TLX4E2dDN
38kVkEwmrnc4uMIcE75nnVCABZoMOSkNQRqS6Mctn50QdpvykmnCBHLQPcOG5IeT
WALHr7qTMa7OR7jECTgDi+uNftN41yItvKienBi0WQTT86YZ+M6EnoyU2kYKQpro
+xEUVMnQaHqxHeIY8JRcEUCJcjAkHfVerOShRXPfX0SE5tY5grWHDDaZg/R//3mH
/y0w/hSKnuXYUrsUOIFHKVDTpyB4UC2XNN/Al+SxWCDvIdl9w8ibX0WI360ATlPS
G/A/1HDF7jKFCPTxR+b+DJilPd4dKd8IQ9eSxpeOE5EAwIFjfmp4rZ7DwwRVgR3M
nJqhJHYvZHJOiDZoeD8M04Ob/RJcQB7KW5zOsycETQddmZ/4nZc1pzpcai+2jZuT
dS+GQH3DNOqkHXMM4V1ehR67bIIWod/mlxlnnwmRH5yas/cbxDONavf3vEr+bUsf
nOrhlYJo/y4KjO2JiRegLPWouBBYLQlqax8TtHde/wso7rZ/T88j2gtKHMHwkGJp
u2AM3tTD+YEZ1OtQM5jgjT8oFEShdY/eQSDeR7GN+szv2nl4BD1J6UbbjySmqvK4
zxjKfmSvY07sgUK5M/a2TKYXe+nNRlSRMdgle9PYp7OMcUGPTToXL49BxIC7O6cU
KzHPTdoi2VQaXGo/rsKi0MoWkgBXZzutHQdO5kFViQYXbJ60Fl9r7W3EvctIcDmB
ilIy/+MboQiIX1/iajAqT2TlfyYIioZk0B0xXw81qAjxfLf+A8Ff15E/6yPLIAyg
D8jeByes/v5PAZGjpbs8D56gCmmLDPvJFOvBHHkR3CNCo7autObSb2eA5m2Ei/kf
uRlu7EFyymXtyspc+65va67ojO0M9uy5I5Oo/oMm27ooBUbEadOimJ4nQduNCx8d
9jP03YlW3BJl/UAwNXUDvxZinO5mvzH06p/k5iCL/lKPbo+9rGzBc0W/OvcbTp1Q
z0sFZ6YHe9jdlzR9mBuk9bxOdT9GvGAqruaDIgKAjRZaHo/BLW3CDDkmW3U3K3VM
bZBTzAnIQmwZsSHbjRjvS9IeNrmRjtNMYWSL9N0QyVrqMNXSVMyYWoXkRgIwB9A4
Dtq3OgqLvhVUha5iyXDFoOyAIXHM7paGG9v9Eqlr2gUhpoe0rx0BBQbVmPFp4+28
onLP9F4sK9l/93JPMU2tK6fhMdW5JjXMaIV1rIFganngU8hKrfGrgjnGvJVX0To3
IXTx1i3LzHfiwQCPWPADiI5ScnuRhid7EIR2xXvdslFxScIcyfE10K93gHQ06DyW
eMAtf9NnwFmaOKY9ZyrBlfqRTqXmk3b3TIIIjY6NGzR6miYZRUyLUzaIjV+Qq72v
vUEyMNdfbfFnLGuV2Fp9cPD+8EzY4/eQq7FO1x9xjwADdTkaa75NfyqbyBe3McPm
c8vOM1zUv6xV3eQsLe94QCjIya2abVs3GrWOx4CWHnWAj6ixUSI33wr2OPNuz4qG
+Mw9lsBYn8HW6ccrWil3H9k7l3vDqkOFPlGC/8AWYgs6cZM4+n6/+rTaYm1DK1Qq
Qa/fyrdVcUlLrSFA/GYRsRkB+b3RRMAWQkXaCgcyh0N4+QOki8iBQQnhyGd9J2u8
fSpo/UWYvc6dFS8KTIOGSG1EeZx0ylmw9SzP4Oz3wDPs/jvXKYdqYLPhpCpRnocE
frSEmlxpK0Q4OEiMlbQydIQ3fmCLTrlQGQ5QyoG7EMBjXzkJFKHJB7/oiuCbCSiE
MhK4jQjHKLBXRKaKHIjby2Eat65FKIvmCSkXn3+4YeruCs8D/5pnHrwyPGOrH9Rq
GmISK58oITDtWKtUtc118kjedeuI/yH8B4rCd6xyK3d1vbAqWkgnDqHduqyy2504
uC8udVVJMFo3Q7BDBpd7FTlJJvTZoR0b5Rbx36lqcMGbWhUWQmrX+kqGFm7PkiNZ
HumAxwv/qtn0n+LKq6T4B82mn6olSCHmPt3YaLjHBTIJgZiMsz12289utckPW+MC
pSODJ5B0GTnKIp0BTvq1HSVcqoTk4GWvM8wtXQMlJtEFW4kninn088iUThc7O8CA
qHyEFl50ZPu5LO+No0bJcUHZg5i2yEnUMoV9s/ZS3JflRpxiGqqzDFzj3dAF76G1
XCNVJtj3w9c5CR/7p1wOiuvCoSGaViWsHmKj0h5iyRHhaZHT3dTuPOul9OE5IKWK
GOQ6Sfc1bHfowLhjm2UzXpVK8EEfVMrn61cEPpKy4Mz58NZtO/qsdZflhLkdz1FY
XjLM5ZlBeLWXJM4ZAtAC/jxA/wE9f+3aB8s9hgz3xBeeHs8osYIvISJwJf0LO2bU
dvwaCmlKx0oTN8Fc9FJCVRljuM/yLCqNmJ8SEh6D4KyTohJGBv6ZwBz/JmajcK+U
U5YtTfF63MshW9rKr5PUBXIDngPHHdQeQCBrhqqDRJG1c8x5Prns3Nc/lMa2/bYA
QidpiTqs8VEt8G6xpRCl3M6fTig6WQoq/O7vkwXObkLg3QWLP0fNGjGPZufHyhcE
9DNn+glm1Ma043wAizRJSsbX43jTBirUpS3eSgKQFw+OuzfO4vyc74Fk2HXLCZdC
Msw5YoBa/utR0Ekw4SBWr536eb7o0+wXBXRF62uV6uaL9z2yQMIoVw0DnqQ+dEso
ieAv9hR917fjj/6OqV/CE0Gc79oD9K3JH2c87u7NOnoatZD/l6VETtngV4CSQfbJ
1vvYTlJ7Dvt1D2AQ2C9qLh3S+RpLbIucYVlLjfLXajy2rNj9tv9ZZCiqn7H97dUi
zX2FVUcvHS77CrE1uRw7V5bzjfTuqvTfD7iiOMJCONQrcMjNopHPrd79rnGbqdd/
jZpxCqNA1ZhMjgFHlFjY4Z8A0Z9CCEE4bGpMS7ZUvBXjdjhS+6m2LKwV0F4yFhmC
Vhm1r/SEUP2t7pwxeohYWB9QSmCnSNYKhfcEVTXjo+9xvm65bMnvFwC3/WuCs81t
p2cgJryL0htGqlJH/2CuqnQ/txwmMyE788tbEF3JWmj1yXiwg7fGYKNDigPOza00
S04TlkAsQiQUodt1CzlP8JS3JIJuqV+eb+081lhN/nrBdKCujK5u4D/YJebPcBGc
EC9eLbyFQcSV4jPz1xoMtPAJEmMBa/49g7a99F6WrX/7Zu1mHVXPtrSy+vJHXEev
PkVPyo3HSfWpCj4kaG85FDSFDw5pyvIpcaZ4ZhsrPwH0rwiL7uGTnwqxUZ0C1NCN
VDTzO+0cKkxe4qbr4e41hBMrD3Jc+8uzdYhUkRe9BaFLuIZusDHzLJCUnh+IwPhb
CKcfu5KuW2rJ/RJA2obis16ILbBvigb4VmqdP5+qIjd+Kqo7ArrWQWcdgipMbW/l
Afegd3aOr877wLaztjExg0HpeHwwDaIGvwk68ZilNmJPSJNTXK2ZiV/l4hLF1rUT
YLVcMV78nF0OPeXK2SFui3dQXpf1SGHsx/eMso1zYDg5zRY3QSmYqHY8nx1axLht
EaeqtkgDZSAucSoS0KN3JcgaheK/e29Qq9L7xYOs2vzeb55Qg0PUbGrTtiwmOboz
cACF5XoFZNApngV4rUwsedou5M2GKLDY9FJAxXqyNX18hJCuPgEasSpuSqAY4Lwu
jkYS5g1Pu22Z6XD/2A59e/SI5kLYH+7BYRqdAajcweVWoT0uevX78ZJtz+Eb5BMk
Up+L289z0K86Bz6yb0YCoroZCaLmXgGdK9M6GW7etQyfmnF3Wi1ELYqp1kvgvMhX
smBzVl+92DxeZMAfJvd8tow7S75i2YHnkRk9/SpmpfgmNXTeVXHBx2wOasXN/CtT
PkcJQYfI+Yx09WOyCTkVKOxCuN/lAj0+0x+Z8pCNKrfDKqS7qm4nhz4iw41K9HaK
qDlnrlPLjUxeoYNkrur/D8VgzQCUGUcHBN8gVHrw1jmDyCtAiawYsPbiMXHhymyR
iPRLvPthCNLTSok3+VNN/ioGjvoOJfwP7SNzjDXPMPmQax0cAEuRHsbtzdV6zub+
/E+dcJYrYJjWouvhYURIlLUTFASEzzYX8iUVFXAIrR3sqUwGBvC02Qe69zBz/div
7MRMTlcOBDz1VwdG7qRXgu6ixEWhv8jkk2NfOctNQUCymwP/ucMVGlk+mD3YnfAz
hA7BZUfphmjuoUTVKTk7pHVdLgRsRF4yUPdXee/HtxprzOF3zSc1rshR7m9y4wLN
EOyA2WBIW7x5NJfgqcXolxj+AImmoz/Lfs/u5bgV/EUjkJD3KjqCWUF5BlYbHkgq
ex7X6Y98IbcvpMO5GOfrg1u4cOJ9Ha6aNq/zPUH83TsdufxveAKMVzQe4p4fCyFw
OvqtjuLICYaWrgpPdKWPw40eWotbCLu3aNk2RgxnoH9Ay0O1ymC+7KVk0GC+Zqc6
2p//OkWGmyJA1zF+bKqZAeBNvJgG9NFNkrdurkFMJZ3hKYOd+OuNWBU5pnXIgYH6
l6FpKmIf4Za5DcMnt788fP8iFVSCn6x6pmlF0Z+3/vhWD3gq3HdMsFwdns5PoDLD
weqUpWkqGuqu0WDq8z4snaKVDbDLA5iT2BimEa+pZbLQJdfn93wpKFTVS9Cryqzb
JS22HC+WeOzGMElxzD3EvQFV/ZgSutLAhlVTWd5bbBjgQMu2U2FXPlMMc5bMYesx
5zf4eomP1naEa049XudzTY0iDjP8cE80enQ13WMUK/PK0H0seGIukrLjrOB64lCR
WjRr89gRgcabvVNqXYkL44ZbP5E9NJzQ6j1nBVF+2lcdtFrAb11nux13xXF/P6k4
tmu0u/y7ZwW+/SEWkBBbebBX4ESDkwpr0w6vi+EdGZ8qQhaJ27V2nkTVZNY6+q8b
r/KIwQt3f4ydsc0qmBntBtxtNc4hHnRzl8tRJV8P7qKw0JrWCFMj9SAF8VyxFmqQ
w0BYbLY4Ye4cufINH5n3NUyGfSLpSx5t8f0ggBDn/ZdgrcOx6pa+RHn4pPtHYrQ1
dzZAx0M1bp/HrxW4Ycw+tmuOkL6PETaKYS6coyzqhN4mFEOSHnyZHwvEZHmEU4hC
Qv72WwesQ/LGiVYYxwI9MoCrCNXDMRRkdhXXyFeFXU4+scFQwwCBGCCCii7QfcQq
bH87hkXcw0zt0gH5f+ybf9u/y0Kj5MjENMkKmX230k0klrkh5D0rPvSpPS0gETT2
iWLullDc93h74F+Uz4CCPDWSGfcQntRojk8NISL2rIyfmyWAnU3EDfoh4u+FOIRL
ofJfUdhnV1bYjF9IMFEZ5Ssli5Zee6TqY2qkVGhjHeqiqCE+4UMKBcpuwTZvC6T2
akYLT7jwAhPEOZyP25eL7ZzlB96NF6tK4kzlaNSRfPiuynHkelJV2Co3/tmNmW5/
yAE9Fbv1oZ4SpDR5dbTa3fhzdXW/83pZcd47jJWaMB1gHLEegn04E28OJ4Llmd5u
91dYQX4RABW8Qsx8+9Bb6lFjw2gEfBCBWiyWODWNM362NhtX1CbWXjs1cnZGb0g0
u6FDypWNuoJcEjnlw8YcMxCxxu3XvPIC30s+NZAVqGYvT5Yh3EXwJPtB49+qs+xx
cT6PJrkGq79TZcepPfIlmoC29P33l023CjCArFDp+HFUw8ZoNFI/Bb1CCQAtyzTb
ohlv8OmhLvBG4E1JziZnoUEdC7ILVSZl1/6IH3MJWsgE6lbmTL4jl4usc2r0qydN
sDO3hgx9rLTvozbz0S99DThiprkHwISDF7W5wbJsoZn++g1hL2CKKpJLGVPdmsNF
PQe0nvhv/5GPFd3m3Rj7MNGsfFtGUKSe57BNpM49YFaYuAZ6/pS3Jle3lm9JXFfx
9KVOsc+C3dayRwv8kdyA+IPQy17l6WK6TqNa2AMNtm9PnVzK5IdDPz+FgKfFn74W
bw3PF9UQCgxE7RZHylE1tNFKqZ612QvGEYxwZ/qm4JYGmoVxVwcZsdAS6CkeYgYL
ex7+l0JhppcDhNEOz7gcXoNxn4Zo7sqbYHoNkyB9JTn2VebbBRNvDPuhkK3kZl7w
lSzWs7qugCgFU+o5139SnOJfsW8i8gonbvyXc9e8HvzbMoFHOUKR7WsNYIupIXGP
JpRiilyWKqxny9P/QKbzIctN0lJZjsLAZyjMpd70Kj6z5lyLNKORr2TPhVKkTJGy
yIC8npAvSKePkptrfSTMLR2C/iDcgxlXkxDr6E33vWVC7rCrPmKzNeDxvkC3Y4oE
k2SaxSMDRqRQuGt7kbmpatdQfwiQV4tHlKU3WEV2iwre4ncMOMy7BAYMmaA1tqcq
PI9QFReRABoFPW6DPHU5gYSL1vNdKGK787c6uXz7TyZEIoAUr50PMv18a6m0Bttg
+G7iGhZjajxD4P3cE9p94iSf94v3AF9xz+uggRY3OltUcTfSXD7aC4xmNYIkt0XP
/BoOBJ43LDcemF5TeePgJQ96GgoDlS8Ws2nNJuq1TXOxcZWfkJsYmMDZnYgQOZN3
NvYHdvssGqDwbmnbYl4sOW0FDISFHa5J8MHe3qTkGuBUEOD+54/jqdWj9taeVzoj
2lgmzO3uPj8Vtcoe1wgeZOQ57I/RIPSJMnPS+4wfNVqt0dlN5cJnegmGSJyH8A9z
ApRmcvd0EXPDOykBo+8toPZAztqAc4V38ot9wR+w+e23IGbTd4IDw61ycnhZUQzW
gdQ8HqUMEASTfxU55qRrbWFrIwCuCVBXZWXZd10s8ucoNWRfKH5sC0ZDEvFUqkK1
5+6fqKgn1fUXtNkXUnZCwEVB8WGJF/heeFJOZjxCf3xAHsuFT3llPHA+LEMIqXeV
52wWLhvPimiHDeVjFQHMuax80V/oPS0dWlHOwkNNMYCVeJSwNdzJGWJKa6kfzOx0
GFmGywrZKOkDfeFGfWLCZ52wt3UOwAhFAchwlSKUTe75RMOQ7NLnpkJEJcl3SAwi
WlmX2mzoKYat36gwM6JnULq/unVyfb5h02MnvNSe+baij2K+zSMzs4TBwzufdYdg
MTX3BpKwJcYhWg6L9TTdqGLDudd73oDnypNfhKXUWITW3v4qE7Mmxf6I79YcKToy
BFB3deb8B8JZoi0URpwQjuoXQtCb7PKF+Fof/beZDsb40kgL5CngpObJL3yLnvHn
CC79bIJB54QuDDwYBNW3HrCYH8MQWvpzEDMjayNIZnyqNaR9AaG1x45m5PzJlESL
gfZvGEGjHR7xRpoC2cz4UNUeoHW5yzNOQk0U1+v7tKlnmConEeJYxxqy8A5T11aX
hMggT5536ebhqv2F6EsMFpR3XzQR5L9uAFxpQGxxlK6K3uUMJqoYH5NAjp/9HUB7
BNr4bn2u1bobK3+wTA2i8oEyRZf2KhgIXWZw+zil6Z+lkVVbwbzrKzu6ma67CiQ0
ypnA6aNfTDmpZaN6nlQj/jgO0mT7pGef2iwb+mo9LZ+4ZD/jfGNHFoFjMJ3Q9Bb9
dcXvTfJWEB21wsZa5SnYt6Xu5l7ukPjv62DXRHlOKZP0qiZm+/dk/nXzhcPVlpkT
TWfqiQgKe5cqNicwMqQ8O1Zwo8vMlwI2oZfr/i3/hQnMrPQ6MlO3BRT9KUG/ZNfc
nO/kXuaeovMRHnXmlIMRbcsp4oDBAxQ58xs2e7D2QPTuIim6e+bIXrMlTKuVRzuK
tfe/VwITpeHlbtYn+P4Fy4Yea7KqMEPwyi5uFpPoW/gAQnI2Xa2+CU7HJ96+0YEp
uk182pe2cB0Z7ppHRRe3JcsAcw9u2JrwwogMsVuLIj0KR/n63jYW6EJ7I8JPRQ3G
jZtnEtWZVAKeFSfJz7Kh1EXBYUx2qych2YAo+kvNV+Hv/qgtymSwaU+6f+dNwBkA
ocAyW5mtf2CjS0wste8oUPzzdmX7OzMex2kXYY7WYb6V2tEiBnTnXNWLo2KyZx3G
6wU8ub6mJEl408ycQx+qkP8qzhjsD6AF7RsqBvqGm+Q67lRs7VfM9GoKFDjpVtwf
UKxrCz0ouqoRl4Rg9ierxLTAQNMAx3WqghBm1o8lV7qHGottLkI91g1dAJ+Sma1s
tGzUpUOYINnDcBFBgByuHqsgKQ/Ish72ROAX+2H5AOVEA7Nfv2GDRDP+sAVL1PqV
AyCOKvR/bWWgq5Zp13vFQwSppl2PDat6kxAHrRZI+N67bI+LonW+5cKZhrJthaLX
/uAGUNAvTaz6y3pJWeXg2wOQcybp1cHcqj443aZtYGnqRqD3WA78zQMTE45MEdBp
FmLYw3D6IBmYz/qztlGdDmXEk/IdLRJCbuBiCSJgRXqeyWUfykmQdo/GgdrSWn/G
JJkERhDyE0PXJ/zPPw8dyCdyNtvWBn22+ykgCv+wwxl4bdtPVVojG3ug/9kq4btp
nXKpgDfFUtdEK8CuTKh8OWkyRMdGIaIHTd/yY3NQqnX3Y6gpfXrmtAFs3/1E9ock
OdH3oW5Mhr/8C+PI5Xy8ZWdbA4kWe3J935Ap4Ap17oPMlfO4F8vdjeA5m9lPClhZ
Opqw3oWrzEOUeEE1T3S4lJcCJ8EUAgxTW8AioE8GRhhAVPzrfIwybnt7DXrZh8Bn
ZgafmmXfUveuJy9CCgLxH1EXAzMuv9mLBHZN3FWEjP5rPGZr+noxv7ptaGPN6ALX
V1bNKsFqTMcASBVLB3JK7FH1CH4E5/KhbALrhZgiHutAdvBT8NP3IibOZGDhMNAv
EGfkrRKPDYLGhWEew4tRSi4s0V9GMgbrpSxzEG08ZCP4OwlcPGSn29nhtyDuZ8/1
fKzDOG8OJUYWEwvf7K3xWWpxmwsqI4Dw1tVHbCU5SaPllS/wLbix4Qlxel2d/EIy
U+xNegj5cnccQONCb9YL9uwVb5megQ8+OsIq/WOV4B9LIJREHKNYieT52J3ubaVR
7XnDeAb7EW9XvZgbyYy/vCsm6fMill2MFlGBtCVVas2kNGNEq8TjM0fHYndEr4fV
jJvmk407DRQqobzUUNg17IUPg4/W4wOWbvrVlEaxiK/SzVcj6ht+Czoxz0YEvg0f
kel5xxhUzblgLHtOE+wXZZOFQs0XJs2+MUWIwJiTrsmJ2qSEb7hppqvus7Kn7xzE
a/MMU57dMG0P2Vh0XEbYbUHVR8vYVxqZtkwsibXgBNjHFUyWkpTXvIu2hzcOeppF
gCiat7+UQxAKNjZKlhkpWpnhyHu4XljGMwAkMc+C+ZtWNjhPZpYajaKqyHwr6hH4
ngJO5x9nteQ0uv6dXLYA1IaNkH7r4Ra4pkrPNEiv03Cm5kBU/tsdzotEMqPD7Clv
HQOLHcGIHEsaiAMjimqu33cDSXgAdh2aTK53miZ2CH8kzXXKJwfWkv9U/DYOIbSR
kulsAdvNpFTf5CO1OyvfmVYObeVyVQILZcikQOrC7gZ6zrFk3d/k32HIKTfUYCt5
p89Z+s7Bf9K/4ML7OXw/4vtI4u8OZTkVvkeqrXm0mvU4dI05XiySCVCB4h7PyAY8
CLgdyR4ahypXCiYKi9g0MiSHhCNXsezk+s/xzN70BJNpim45IAjCRxgMtqaJjVYC
fg2PGGTpJnaM4AIXfj194+rIzoljuK1tQkEFqu0uodRw3c0dChyrEOA9VUOZ2+ra
AMRMVjrl3KdDtoYlY6is02riPs/g4fMeijUFg8DkZF6PzWMCWxTKwOZ0WA9GQSYV
aQ22LPvt50eCNtLt1VdFThcHmmENW/8H19OKYPvunldlTfLXcJJqjoOpnGEAJiqk
aYRnI+zwyy/4sMzM/cyDDtqMBTO5mz4NAnq8FbrYH557PNviRq1LGpIORig3MuyX
O0IZ8c/R8ssa13k3N47/mI8rdI00D2wkxQ8zhYcgZR4ey6UCGGdIhtNflY2ppHZx
L5UdUBl+JhZ/F3ObJYvPjPMPz5RXZjaDnQHgcleNq1NiIaEPAJCV2o5XLiezOJoP
aJXnIpane61qOs2GU3yOqsqOGxJb0hpv/yLtHNvwZXjKwp9jnIePQTjJGFn7xQEz
sqr6ZT0SlUbfshjgUeXgZt9EPM3KMoPPExrKvdwPDWPdv04P/aMm/e00v2o7AUrI
y3f05oQCIAsfQj9iI7+3Np2vjJFZ6nZnkPH2hE1U+qYzNpZLcJMoRlTczRS6snuO
+AvM6ATg/I96j5pmBAJsYTVOhbB/yS7K/cGrMpFQQFlGx9e5/f2NmIP6IejaPXK8
qfs4/PGx73O6itdxWhydNWKML9lybxoAWTr1TLlFWHheNGra0D6Oc4fnIbmRpRXW
YHennqMu0W5hdqYJFHzw/Uh0eyQ0IFOE6SJmL5IhnNDDaN3019PeZiYEWmu5OiG/
O9jiNUvHrlpNN/KYEA/0HVsQhZLwGLr65RE3fAcXbee0oX/B2/ga9TaRkLG3V4Hz
xctq54TpAtEL9UO0Iqw5WJGieXdW+3RrviqLAvC9c+8Dro5ckhMNActY8Jzdo6S3
UsPXTBGHFeIuoy/C63g+nGXQZcVDnHgD9vSY7kgxErppy7yfnP5bqQcbVgDRb0ro
NVglIRpeiu0/ayn9dLxi3y/+NhdY2esyJy+TxzTztFuNtdPbCn9xOQDXSlAp1iFE
cDjoAc8zvqtop+UgGfMNf4x8YJk1I0xDOdoOgn/aQ18dmGUQ9UAR4mfELnTmSHKK
jfktVLb7gNAm3YfrVLywV1Yj9hs1xPMDf0Dz/GYvnjXVlIyr339b/IA5SYX7eXVo
14ezwVMkFTSg0lklQOelncrxTjx7SFde89Zec3Fk9OB2D4gPe99PX4/ChX72Pzqw
BWQX0Qlp6zeKj8ow8oCXe0F1WtbWNmnm0/MXbhGTCAnKV7eKqRre1n1axP4ChLNG
vaEzLuNPiTbzJ0trPrBVQM2lRTAVvyGvdpIpodktMgT/46HVOdwk/iKNzTe2xWhK
XjkVAAWVHUaWgL+47BntHtYVcNJJXexqPByj5iHE++Oh/BeqYCKGG4Md6ejIkuIM
/Kxdd6n22akcknnVSTQFhpZta9j57sKRFBp7OAEQ9QhtZlJpVHOcCkgpARp/7s1r
6QRYnRqgGcdTuUwII6isnuw99cHu/P8ps9JpAYmFStcYlUf65XhvtIBI9FLw6TAr
XlqvxlaCdtacD596PLI333+CfBIkAQorGSgBjofZPDSrR3CkgbY8HO+bhRmrFO4F
FxPY/bgxpuhODsuTbGhVBaaMT3Jo7ha7VgxDLbV8KLko0l6nvaGadyeLB81KsBNr
a/c65wecinn8+dYUV+TKCQc2LndGmNtVWaZjw5r5txUKdRnk3xpHAoN8CIKI3JpQ
2dSOge3v1WmTrUjsUuLBEmhK9rYAKj+QTm+v0Zf/UrLlYuFKP0jVw8ddRhjNgBop
8I31tnrr0DIuvSZVZEySUrBa2Bdqgv5X6nqzBZ+PnzmYm0FvwpCzDaiWSe/VXap3
izhXPVCKsrJIIUJ/U2hsO7xoinY+s0PvGAHT0zIfknbPoB9C6YOF0fkJihszyQZ5
y/nF0wawpMbgXXM9SlrzjpI6daCY2XD2wMo57oxAZJ4wNRly329KUGXv0BXnex7e
G9A6VVyFkSnEm6LnImy0k/jUcYMpPYnz1yuV9HXUrAft4uuQzu8ZzRj4XQYSV9Lt
vEZQvNQBAtKtxWzdhb7ZYkp9034jWhRRk+dsh+6LVHR9/kOGyU6T8ISwJpqwr0zi
vXqQU1SIt33ESdRHUXe8ja03kVbtYCjSvj+afRksSCiLU4Edwz52Bndt2bYENfQg
18Pzz+KtZ4Rp38CnfK7LvyS/W1+HzSbB+k3gl5B5SU8/C/iJTsXNxmnXVLz4QczV
Q+p+fkL9+lE323DC3LUqE3qG2+0q/beXckXTuuFLdi/wdwm0YOoi0HWZMZHEJpSm
PgfUp94TZdZBplUTcXSXgLHQEsTtRYqdVTBUAiWi3ntAMQB3mEA3/MggAP0xrXid
o0uyKqQNXBuykmr+jRWNeW4iDdO0iDFn3W9kjSRkemY4YMwJ3dVDFMrG+RpiiwTf
7x+2bRAZdDDPOYLZqGTqs4VdtVFfZ7LgJU1CbXA9Me3/zHLlHc33CzsTcNzEeozD
e663c1gykjjXCyA5FeBRcOYCRi32XvrtQh83jszQf9zx0XqnZOv5+Iorf8WIrLtk
0zZ2zBGlCP8VrJ63YjgB3lA8uBbTvmc7J+UALzJCnqpmha4Jpjxu2WQ2+DljLyg/
/SmapPkNZIWDDu0AaSlAPvws5VVAZjeTHMSLNKqVQJL9JGiZ+qS2lD+yYlvOfr6S
jLN+QjISDpUgI951U+/FTtZTmP32HwkdOeYfv4VYIbO9DYAEkKLX40bM5Uwt7pDp
sWy4lSGq1gNFcilN6Io6JERpJRjJkH4Nl2NH635meRRd6cdh+qrnE3uYJqIGH4H2
3y3zypiUWMXVlXmicUFHlsAXp88KL/HrfoO61fiVOvhcCn1j1OBS/8isAdLB/flp
DtYponDXc19cTytgsPGNIpzpNEWWaGLRwZaVR2zV9/qGcg6ogfMnnRSMKLUX8nA6
tEY05i7bruCUokZpt1P/3vZfIlHw6j03Td3RC8r2dQSY9zWFQ7nF9tOy7qUEuPVX
ii/oP64cS2EQ5HSws5Jx3b2Xo0DQbGOCvwo1EERo4Boz6X1yDOtoY0t+MPrj3S+U
TGLshVSVGjKrT+pQlT/+oe1eEnqrb1AebVdiW8whRDzu6IUHM1a7qs7ZsyrIwLgN
4OMGe4SfEjLIkk8iOeKIHhzD1GsZMAeuCglAkwU9iHYi5du0eiX8IBJct2lk4wwV
l/JAG4EN/zpMoSNf+1PY9sZBG89QPdOHUHkqtn5B7xM9nrMHfQyNrSncQNGvRqMu
oZ0CnJ8BuvGzlWRksL26wE34z48J5WMqP+cnCK1b0twCD4uAHSRYAuzcl26vC8b+
vUrH+u28x1IeoTW4YOQ/y+Ss4LouH/OJHF843VWg+YFfVoFtAbDNpXRnZNjP0xQr
RVEkF+DD6E34zjNC4bDxvIV9WSKOohdkQ/WbbapIydlphJ3AcZCZsbd6y9W2/uwW
giv/5saWU05gL6ZtoNCS+7yeQgJeAD2QLZc+G4Ip4zLWqjvodvK5g4id4qAETRJP
8UEktGWMQ46AUnHC3BLfBNYfaGZ5zPNu1spzCU5RrBod1Khea/GAmLq/eDt1qDLg
+jiTZJCWl/YYvhLjvNV1l4glmZq3iKA3xYoLKE+IXBGxCgodVkwuack6nQZuKw5u
1TvqEWFpPYjgUUfftjnt1DwaFHCqEyrH8b1DUdlyQCjbuA895s4oLKdefUZ87Tyz
DwYHpj4Qj47Xtq54g/9vyAGtZtolrgOSjc4CTED0tY6YxfFRqo0/2tOALA2+HG+3
UTVzbeH8UZLwXME4ufPtf5jwcLvtoZGbKxC/2gLFGYJeZ/Qg40cWnZu78k74L+lV
JWirJ7OmbjX2sinK2hoJr47a0JxWn+8/QXTiX/3UYFV7/X85bPTW0i2iwJmD7z+g
DgpAHi2mQbdvXL4KJ1Ymfelpi04pb3UjwJlq2JhJyK0izcEk9ZDowVwyLlJhPh6E
JA6hMYEJbqctCL9jAjzYmKxIjE/SZwk4+WS+99dn7yM8PXEX2CpNaW9oeQqytp4R
lcG8EN+teh751ABFfEbXfrow34LZuESGsG8R9Q6mRzGgH0xs/zQnYC8bePhuRDlU
1ecVxvdIfMGE4EuTDV1hftEbY7pk7W6DOeFjY0I3WVsH27S4V0RkzRRWR76Qj9nD
cDIhgKQIOEF5MGr1d/IJ92nH1SkjS4OfdDu5pcYtNhWTiw6jt9gdt0mCN33vk+KS
YKc5Ih6GPudQuLBxfrbC4anJk2Npm/LTVk7llCXm9Af6/71fnN6/6+32xiWX+AYD
LQ1S7dLgYWOf/VL/2vYLSwbCOqIMgRD5i6dV33f+vbIQ0EER9V0+EXJMSuiMt7QZ
Nem0ml0qCCD1BJCjo/f4PkfjDW9lmCI4qyAGwlk4E816U3LkzKMehxSc5uPBeJ7/
buHyYeujqlgF37meoa0whbp81IoRNTfIL139Sq+8V5+v+A8IhgXZw7gF/h5LSUu2
KC3q/ZwBUJtZJXCMNHzJ+DPsZfxw6Rd0EDggJcnVahu1CeOEv55KDbQ2Zx+7lurn
wRF2pyISiLUHfuME++157xUjYj95fdr6ccl0UbqPRWJ6kvfI7JZuLeBmHjeRUlCn
FyXYljbmCYaUYS0p0atausxjWgGsbI9wsbhbUqbzdmqhteVUj3DczDbMkHOWq+EW
V85tZ8tvQO2+y3Qjf+v4u/vj1VKeuJ69iDLOMmXdguQM4GYzcxXk75CFPBmnIjLw
QIuHCA0lm9Y/drq9FXhD7CqmHQPBIOVik4H/il7IFfsyzAhwcnE1nj9OfBcgY1/p
bGI1/oHaHvHzRilcLrfXNogjR68qPofbhhWd0U68iaAncQpSSwPAVDd3vatrBwg6
PbHeyiursMofQ7taMMWRlL74qmlEFmj8P5I+S39tIf2T+yHr7owj4JEtOCJKWwRy
oYVjUirBGYkeOJEbgLJ4mn5JCJzY7dqJDLg4XLYXn1GNHI/Jfc0o+WATb1JthvY0
Ize29GXEmh6sk9JpuHYLbFtN1YvqxaxcMxIhi/dk1728W0ZO88Iw0H0qxYmPcDre
32A/IcSh06l3qyEOl554lby/Ei40Wia+ia9DM89/Q70Vtdc90y3hOit3kqFexCfC
fGb/sxhPkkdZTwuU5culm8ZcRKY1yZLNPWyQzZ00Qk3TbomTjqGzJvTBiQp0b7pF
PS9yCSGVI+pf2CXSxCzthB1eVlE1F4yX02mBrpe+kNX8aACjpPwLLfikBvx5vG9o
WPClBwwYpV0+CjBn13rvJmU1kSnWupVzH/EsY349wf1cUFeuV7tMn6gKodTf/UPP
ukNwMcClFgvCex6UpkTdVuDNQjmbLL3bXIWTsNS8BkJi1uMQtWEekbURMWgvlGgZ
+BTi6JUjg55QBNZLg5kd+D5zvw/lAAC6EiLeKuZqvQYxggAqoHgTPaZmBP9/s/an
6iussneOJtmEeqNhii8fUNN+kQmfWVuvGmv5jgqxrW7OKwCPMXy7K2/KA3uyYrIj
xlKii4iEXvbIeXSLr1uZlIx0raSwMgRrU4lDO2SyOL2ftMAPV0eJAEz3Wgm1hnGn
qkQvi2AACBEA1wjSZ5YgA3TV/N7Xl/enSRXaOvMUrovIrYsaKY4iYFgCdmdJDST7
EvapDbajGZ+q5vpZssRzJm5NrRpRcb+WfCnUl7tQjoaizpKV78d5u4xWmFshN009
kypDreIcZYC/V04Uf+BwkivHhb4u+hTEmN7gJopKxqA78REcPDOUDR0dBmmjXbx3
Si1HxKZ6qwn+eMjjDWrepFyDUlX07bFtu9CeyRvU9A/95BKxUUlltM23LoMuYQg5
xeoEfS/uM8BdbP0hewyr5b1KOv8waBsjBAN7vhk5E32qnLOBLyDoM4y3b9O/AF8A
kKNjM5U7M4fQZtbbb1IPKCMa4DtSvdAOYCJsb1gxfFRZESQd7BewaSfTligzgQCA
Gz1wpaM+f6KCITRhEEjoEUV21bHAXmBjvEMhUsZY7UJq+fx/U4oWKLRzPa1/IMc/
QMgLQBpuKCFYs7g8HTYn+/mGi3aD/5dNNxhyHxcCTEF5CSGZ3eXWl8yw8i+M5yu6
wbdhm9a/lHzdDQ9EIC/N6SB6n0Nq/bm84G0skxTubE6KtdVPxm2m9ZA5ODpsfZ6m
26ZWf26rD95DtJk8+MT70HXxZUUS5UsOqIOzlwWE+71GxQJ5Y6mST3yUx8ukcpMe
`pragma protect end_protected

// Copyright (C) 2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
// ALTERA_TIMESTAMP:Tue Oct 25 01:47:30 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
UyDWjImlKUKgAlKK1r4Bxc3yTlOf4KXNuipeD/fWT8eceRMJSh+NRAEATsCIBjw8
qptgeE91cX3IjvPfvaqvjchAwvPa5yAbAZlc3GGSdkJl+VJvkLGbac+Rudsw2SZK
8j7AuIXnugpdTqqXGd+BEENib1jvBQLh2U/wM2BuYxk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 15696)
yaZwzPTTFmm7drfLgPxlcQU6tXvKVL/1kW1L+4mK/ro+SMVRnPrlpUzdbAGXTFO5
9U5EEOJrjZ/JiJet+GrKpPlZrLDH2Wa5bkkTWti5lHIHNytoYNrzzvp31G0SIfRX
ntMj8t+69z65HbiYJSHjJozpE+t4nVtXi4ZA3nklMQNF2iJ8xc+QML46W/Gc3n8T
dM8K0zciURMqOqCCswd6slfNkHesk8l19eZkCo/GMyQ/AWfiLFbnoXCe29A3rCDX
wOaaO5cymIfcXIUJG1hW3575YgQKN1Nc7WraRQjs9yUWvRk6CETmBANYccISRMxO
+4JFk13f4wu7BjXOLXvLwRzbghGigoSKqfc7S9h8OdNDC59LjmDkMt2ueH20Dh04
YNqoidjc53mmfeP/z1oNCYZT6NvNkLZSS3LdswqlbUcANGhat+5l6OZd2Jt5+Sju
fSgr9SRPOR0pVjqALLeUm+siWKR6pUjwGjWt898508dskG2U4UxbFhAirdC0gvTq
QJ3CYs0Rh/MEumVElF6dPe0v4nxKogwmKMtPm1UIiNQZbh8HtY+5a0brjqE6bom6
rRL66GDlAqAa8CRtJ5bRHpuljOum9mx7l5pEwmmUK3/eX40iOV/1TsXvsg8IxA1x
bQiRwbU48PQqSc3tc+1hbyMxOHrue8KpozVz0/KbVOig1opA9zWC+5f2/zP8YRIv
maSUe8g6kQSDdaKaXa2PJ3TaDot2f2vq12mPNGqxLlIeUILL3l1DjgN3JGw90Pv3
7Iz87mSiJ/850jbwfX7BKbQeE9othQ8CG1Bc61S5EMwKeLtRs1CAPa0wTjOu3jPB
LXChaFk3IgJXF2lp9s8BCyrknfJhrlMab/zgBjb7x8QUeJdOsrjbQXKU9ryDooGj
iRXE2shqx87yPjyX+bJi0KtrxWWUl+0s1Q+5NC/o1PFhOODHmW+/3CuibkK2CLIv
3fOK58PQusGPewwNT0L/icNzEVxIF734n0Zg7pPwR1u8iL32znD9pzHLXrlKoMMg
cXPUdiJs5/iNJkYcjz3K4xrTKEwYxLfxRqQn9yjUGTKGveGhScaq9tVUXdkGhAW6
dRQRnE0d6d6L0rvjz5xBANBBiNPAC1h8RJQ6pH3p9j3EbVnAGVv1zI3R3jWMa8fK
xic4uRqdMECSLpYm+Kfi+TwcjyuBVMmCjhY9icHEZr6xER/p1v+O2Jjv+H4GqCyD
75r9fh3HlG1o5JI8jI9FXSX9zDiXtjNDyMyMPUrfqLUGNjqAhwazjJuaRPslsmbE
7EKSx1roHvFxCRu0Aib4hTLG4MDb/wMjh+DDtAaRQDU0hgV1fPIXzfyuRhr2YQuL
nkTTZT+mRIVO7Ki6ZI9pXsXR91EvskRw2WQ7ShmsLtmY0Mn9k1OJ7/+rvkOkv5IU
TmS40e/QIqqzzNFCKsFEePh5ETPkV/Iy9giPCoS6fMPQYUL1NZHDHh3ex529icd9
SzSFad3dMzrxK0Y7KP01HJstbidqAcQh83uBeqb4bO9KL/y/m1bWuLE/mXQq6HPD
ZMEtlqEKb3KvHVqeus8FgLsZjFc8MfZA5NZtbf/JoqGb3RBhUxYH9WeQ5rm1BK2W
45nX1E5LioQhaZfZ+ndeEWZ+VBJqmVUTIAEeK2MZAHmTqDpPhVPkTaaEZMU0RJo3
S0VuG49XQGUuGF2NeG7lsGAEOJ5APqd8VJTTkxfgDu/MWoUy6L5WDsuMOp23uSFA
3vMOf4kd0OhruEDKOx6Q4M6nHSBXR8fS973lHKb1mbn180yWHfEWNvXmYZITq4hO
Wc9D8WgjbLPatmu03u99ZvoX4fMljsU/MG4jQPOjjCMiRv1eJpiYaHMZAmWHSaec
oFFFxXAxOyMVUnRi/eKCViH8whHb7uKJ4l0VPdtrAF9Hm0ty6FHn+UAWUD/RBs4g
NyKUVQuh/+LoRPx8/zbd8KTEiG+z8D8b6kDPsL91JAbhaF3oTBx4mUrwQ8RcN+pj
7dObJCd1XO183kTpqfnsAV6W87Depj4UcI8EOQxLa7kFu+ZikJQP8d26WH1rnHcp
bVwJvqGHkGGJ6fT82B/m/5JKXo7ZUet1rFT4bq+aqvVrtv9m3ivfRiQ+hhXOEDHV
kgX/2gHrwIIGeaLNWJpAzlGjsUr62eS8W0Y4cO/unrOekGKcsF4O9jaHs6I49MGh
bpPxeeEyumSFYcYvbwi+NQu8zPDyKzcMwwiSuSz1cYw5e4ekGFhVb3JB5AIBdihA
yA+5ZiDlXIxNkmMEjiptT02qRvQWS4dBqtSInQSwMnwdJeMhKaJ66JYjwhZgn4Oh
6x9OMRUo/cSc9mjVqJUquLLKbTDXIL7ym53fLgN7q59WVoLJ19VgQUgI7EHK7pHU
cgB9gvD7XIkQECtVqaY0vvKh6ZQUbKDtAOzBuB8s42m0c4TwC4wUOywDR4lZEPSg
dlgalYPpU9YGcGMM9d1aUiROm81oikrTUuGrZUiLSZW7h06EDIVAPz2muVniCuhr
L1pyc8RvB8GTJoLEtDbhxxsxWL49fBMxKdZ0o9wUzYlB5KAXkGyH9Ix37C60ILfi
a5rBidzhemNDAWH9GGYVSGt3XUo/FUSYR8m9zudI/QainqhvViwgDJZIzV0qu8fZ
4WocRUXpQvlrqs4yuEsLZBYWsNvTT74CyJtXgAkksZBczfisdFBmgtbLIMpi9gIi
bTa8tvtd3SSN2WiW41v6uE5u0tNwNJXfsGU2TNRDLxPdLEHtlHT0i55qzDA3qKon
V0olC2/HTsdyDZwxG5FhRhrjioGKhC7DT1tk+8sYfPUl0p17kgqwRtUc52rN4k5N
JgFdtR/9lFrLBlLJ9EcFPQLxtHZ2ics//YZOnWCv8Na9CIFClDDGkGOtsKKn3JlO
GShaapYddyAOS/8jhjqGVBL8KdqPeg3t9jssVhVkc/bDzM2jxeaJgoRI2Wuzzlj8
AEKlRSWIDw6SvZPOydqssu+a9O9UfgPTpgvsiiJrlJ6L2PakYa71tUuz2KEYkzjv
Mc+zIIhDrQJrcZLvJior68/gsVfzVNg6hc4IXsKp2TaJS2KkvH4ySyP90dXE2GGi
UoSqcoIJlnaJcIiK4AmDj543vdn58dzKBxcE/OoUmBE4RsJPrKNmRis+Q5iz8jNt
lu1+1W0BYtrO2Ft2M9GYeu45idnBrsMXdQ4ZVi1JpXBOR85EzCOeyN+6TyrjD99q
4tELv2ERe8TZQnFlBk7LePdIL0/J3ks901XsO0WcdwdBMNQoXnQZ4oQJF/0qSZej
VtsXx9SxbzzAZlxMEhlU0FbVbWUrhJWUAR51SSpFaSnFt7b6ZAflD+07F2oY1aw4
3IJ89c50bNQMUu+y+XoNO7dUPDcknd82PIXuZ/AgfgUIkXnbhgqsMfcmjQvGX0hN
LfjakO+/EhvAcXHliman8lQcjnW/9VT4ZOXprTYW565VRJaWnAt9ZQwCtSPGMDRM
yQNS0iFVfJvkhpQsEAf0hKmyt7WE6tsD+Fkb4VxS7wcgWU41T3r1x/UqJIFxfMTC
PdVilEeksfMS7UjKPCc3wmfdYDFaBr3eKVxJxbifgIDoXkhQyMg6zsGnT8TUvKKJ
RqGhsAgJAsYMFLwsD1peae4xtV550IGr9qooQCXm+Z4E8/uSNYJPZI60iMzkuDZ6
iDxcKOAXI0VVjsVlipOBepvjfdKDVeFbz5MU3YPSTZcijU3b7gxK8QYLPotKV6rk
Dy6sOtiKUmtOfB4u/7TssTNK77mbiurhzDXwAj/BWcSgS9/xaYEwOhs3yBx9oOtk
xjFgpP1YkYrZgsWzwXyDzPQ67fxMxFVheB5awJ6dQC8gYHe4rxCA1p/M5hjCGzwl
p9YJY9Z+ZdRmjkI66gTd8kti5RKAm5JVuQ6BVaA4ffXVZUwnDlAAtq1isYz1Qz2p
Wb1MP6UdWfy+oNFlS/BCjmrHyDVgXuLBNpql/2vCmR4pmSJNacGNNvLrabxFnubr
dH2G4SuRzxwuQpCUWlIzpQIPSB4CaZ4mAXrdVzx1MloYFrFvyMBCfNo1xJFhsmnO
DlOPAxJt3OBctpH8dAlLSMhLw1qyNT3uDvhaAgiWcpwuPnt9fonmA0z2O6lllG66
aFLFTX+Y48trp/5DYS22V56KTXc7EVK5KM6SauBd5pUIBpYRey6TgIE9Yx0KFw+T
sgFj8vOYhUTCKcmut3a90Y31XQDF1VDrEj+KlSicb9MgiR18Fa/MqeAqHfB//luf
T4zFYCe5Rl+logJOEkHUxdgVsnaCD/0oaf2FDMDic5AUm21WtxanbhP0CxKr1CE0
4WgiWlUB6MiF4QI5q2HQ7PHBbO3kaJKnlI7cxvXe0jLgrlDo3nd6hXt0PAOhKSV+
foRUR+W3aobxjNK1ZM+PEBaWxwxMGJAqrgma+nXft7wKwfdbLNU4TpB1j46f2smn
UvKyfYQkx6Q4T7V+gZ5GcMY8sRXO7MZ65BTP2M07SCRztrwiTv1DjLDQ3yODkEnW
QyxhRLWGEexsEeL8DoIZPjsT9EhR5XnwwTj/8fbkeo0D17JDwG4YUGJ+zfo42MUI
lCRH1GngltmZRi1Q20VJReFOmp38nucBMVO0EP/cV7sIsdFRQsoSihePA9fp8dKS
4qOyMx7Co02OsnY7t77qkjkr3JeCSBKATEM1T8XUG586CLVIMA7uAK3Q405X3Gwj
9hmxJDAEZKY7SbL/CSs8uKZ+N82dag93Pq5Rr+VNwM2spG5OwFYow+CYX1aulKN+
k49Qi4Y9/bNNVRtzYBiToOXIw+Mb6urs78EgeneOXEvXvY2h9Vm9q8/M2oFsjlfw
PuvPxwaBcRBl/Yx8IDCmZSuKApynA3W3Q4i3HBAqq/QOuI6LhZ2PtXpzEZx1Ut0C
LDv0U17h4hDvy7vi2JbvDUVR61GEZyqKRp2vK4XNOBCxDqcUHQxeTdRedyGwVNb2
DMKkNHEdCfD5uRM6BMHPN/qspjy7v9uE3E3TkBr6BiArb82Dh/ra88v3wVB2+7jv
31G74OEIiMhdd9pqYEJmFnbknD+5YLGExpTL0BMMAlcP1vDX/lkp5E7USZTL3Ni8
3Eb3Cf1BDgB+ixDSX/Ul3A3hzGmAV92yXDKXK4DBUiqpz7wY+T4uPmQnZliVN6j2
g+7S4mlB4qKy7o2s/Yt9+m5wmkejpSfdh5AieJwbjyTnHaGhfs2mlSTHiqfbE5Ak
2ZY925e+mcUDIqlbVcfwytGYotCwrcNwat7sPaVBRn6YKW6+yaXKpX7GA27Fxw//
mEXFDTHx4V8OkG1hahvmO98+casHqgWXPeDr/jloy7cvT9Vi9OMY/TnSKL1M0E89
rlDKN+nKw1lT8Nd1kFqC31PyfFrgDFC3VMQUYu3z+aYCymhiGZj9i62O4CjI4JlB
Qm9JbrdqLrLjQWVFB7XoisP7SqluGh5eKcyDMvTAGF3OPyw7GV6H2jev9sNGFfEB
9a2JaZU4QV3imuHSTwZev8BG3YWQG79zSKNTcD2qQvZri+arZME746nKzOJUFIEH
li2m+tnp1LisZt2P7mhy/5sQvjYhFGJPX9LL3hNWMGVuV2/r/RWse2P1rmMNT7ev
sqEbUdNf8BwHXybFy1+r4vozJklKUnAA0xU6QgiNjg1T1wrcUxDXAROjqW8ICLQi
DHFic5mpM3a9DSg+9y7Jv97LNSlCNNtUz9xu5vBLepOGVFbqVfdq/71QfIP58M20
7bmKoCYHy642scGu5LgblGdKqWactSdItTxVSpBNK6e84nYpaUhGKxAOzdxyCNS+
Kg48O6zAaDolcCi7otHKox2k09iQ41e6RzTZ9vBKcndmGnzzWhESSUGx2JgUfUdL
q2BU8ewLPf6tV1HkSvyCjdT2dBRsXCswtipIVqXk6V1aSoof5yqSCVYz907lpZyz
1shSDfSPBSOcYnwEsfmu2DkEAX8cofCDFVHx426VtpkrWtpKFTnAfrF6ilF08b6h
rIJ/O557BaJznNTHhatXz/HTewnK04WS47gyyr0XJkrFWHy37soYkngt5Qbh6/ZZ
U+VeWjAbH1YJI0g1xRTPVJ0rN5eQVkIAlSlLVOyyy2FtrjTCgeoopTW61uulAsvd
tS8c8CqTlZ2rZ8QBv6frKK/95AK1vMobPc3/h4djXIYEdZz4LqZgMPodKph5O/V1
yc5IXOyp38HjDnJtvXlHySA6HALtuG2H0iHp8twx8BM3ZTfSc9djbhbRkbszvK3r
971Yaq4CitCd9GUPwaYn9kONdpAsaAjTgWoUHTovaA+o/8geqCGizcdyjhW43e+r
fKcvqsGxe+elsH8PG3yTaDhIa3BjGq5d038yE0SL5YdicbxVIR5wNU6DviofHEIg
liwvzPO6jfMERb5yt+z0vdxkgZmNhdSX4m1TLcAIi4K01q5ra47oEKmtRoMSzFeB
XimZZuyNFdYPB0oK+OvovljdOzbemOSvmBOnUyXNobEZWz3vt98UoiMpaFTf4fQg
TWQK7EqXFam2eOV0fzBDglmjg2GtkWF8ReEOxj4dh+ypos8a27gy7Uoi5YLCVob8
WZlW07I1drJyg0fAZphGYo2I8NSv8jrt5JoU6jW43Gr6JaHfjbC4UsAfnWLFJXmx
6PGzMZnB+eU/THA0XO5VAKF7I6UXDRRfQ1C8WAeT/5IxXdSa6fjO/twlTC/i/6qZ
wXf4fuHGFT9461fFH1Dge8Gw5un0zzM/cW3Iit/j7U5tfnpZIb6wsRQwWVgcrev0
jwnL+GX4Qg4JpQVVD2sGwg9iIBffRgOtUJFMFrg6cFJUocG7hS+Yg6V4yiH0UzBe
ItjD5sAa6hs/IsuZT50cFS83Uj8dvQFpEGDy/2D4C8eArNa9vGVGSWe3AoZcE2UF
szg9QNHFeR8bR+o/uYUDVuRq2ZKjd77ZRqFTZ9f9MgV4snEvhs88Qx30rHsgqlck
8QT8rBUioLmynGXPXbr/WDqwhh/lWlvj+0LuUX3K8TlyZs2e4DufobdlNAun/Yfa
4W+tDlztONCyG7OoFqijsm/f6t6nh1ftf3PmZN6m15K00pi18oy0ViFM/FsQS8Tt
z0R2pPsA2Ag72QB8oytHfC3O/cYd8itqCVvdX1cm0u6n4zhnqPptLKXbqiR4wF9/
SFTKeITXFTS2B291/35UpIqWzud20YQHl4/5toX6SCAi9QjvtieN7wL5hgkMabCt
OcRtyGat7KAlJlyfwbQhkgbGGPmcrsk5rYjHU0HnjDsEMx8cBp42GNNZBvKYdTNi
Eextjrr7mMxIWBpIXUIjTq53mRDxTK2FIKLwa5uZ4wjhJ0+ZYYBXQAFVLpx3ib7b
FszwHek4tNfGH3lYed4T0uR0dVdOP/MPORdJgr8iqiF9bJtSFnEdyPM9yMXPRxSv
bGnZ09pVoa9/tc2VRzfeur4rvrYS1re4/Ml+9vQGn56Xj5t1ArkgSZ0LvqtMdoai
C2UZuofQyI3Jfiatn96MnIR99uXX1KJhZ8J8jlEK7BWimgaGaEv7ku5MJWZVh4sA
8xPGcH7Fn3VDS8O1wa8XkUWTjJWj1EZ89gG5z9yu2bvkvmCYEMRj5NjkCumYhSBr
3+sDcsI7X4FHjaK0bYt+EecHQsSGi2NOrXsVdCi5f1cE4QA6wYt3tXuPNmjAFJcJ
Hk8/bNLmUkYms7f69R7PjLN4RvwfFICKudpGT7n1PQP1luxVBtuAt1M/675QwF81
96pVH3gHP3qwWWypUV57X5EMRCknenvmIimrP43NiYIowUaKqF2x1e95Ci6X9EJ1
G5aya5woTAoTJ8UvwGdJWvS1Yv1wtsINVc/rSBjiWshdThfANxLjF9UZFnmzpSBl
hI5VN7rXy1R2udiUnxaJeyGjpC7aRY4kfTC262Jwse+idVCv178QL5YD3U/d/l7h
Fy4O2EBI3wQr2lwo/WMAgNWlOv55pvXBoGJ24A8vsI7OtYfsLFwy2kJnZllEyXYN
51+ZWBNcO3e4o6sio8xespFfEKZLk3n8odE4LWEgGWO/c9vj3w63Xi8QrfVlmTlf
LYKDezWHmW1kRsn/9VnJHiLclgAmHw0GqJJTEIOikLz+KMk0ReosvCwyK4hoyZBg
D1YH6QwSBIRK5t6Q6Km6lKm9Tdyu+O94rndpYV3jPf6/pafi59yT8iJaFldPlRVd
RwaVHdyAQvA7XugnsPrLnbIAUcZ7Xfeb8QeddQgroxDXG/TWqekh4kIsnD2pw8kv
Hh2DioEiiqTlLtE17+UVL9oKApSIeM+x3fh3hm4iOwI6OgyQswtvDHDOTK5Jl1ld
xavdL0n1U8QkMHAYTuo9qbHKkS6sN6skfSMpZ143y1OvHteQcsjPi1jUvZ5ASQai
R6HmC/kSVNoLtsqOoZ7rMXgvvvFrBHmONCGlonrz4No+rb8Km8+62y3DYjRgfhXi
DbvtkuRakM2uxgNscF0tMWDoVyjIxyg79dDiFkYUThIdj3rQLJCw3D2yuxlcI9GI
PQ30XBi1CuIz8xUHRpmLmItxLdrVWMwtxn6oQFn4uDJDzSYJ168b9nMG3e/c35A0
GDDCEG21GhWX0lct34djSNgZJFcM6wXgwE9PdCBcBzuJNuAiny8IqC2PqgO/U91J
e442/SVhv/J+KkH9XGthhMPejWoQzmEBDeeOnbmpnv0hK3In2rZWUC0H+lYl7IM5
AQTta9a6amF7g7U8rSgFAmkDozau0DiVsTdGhUpq30gNTf/xRfF9kWdfRoO8UDEs
NVd7s7BsLo1WsKUgJelrf1pFKaqfdMQIlNaIjqX/sFVdpwKO3UcA5FrjR9eRa4K6
swMa9N+v8BiaIMjMdAAyr0ljCY6miZi0C01sl2aSwgIV58Tx7bWnadoZmOLzfh3U
8TfB+nuMNPeWuaqVrvsOsmFp+JnKyNLSwkBgUTg9kKZqQRJqpMf0yCkM2UiJKpFq
A0ZZ9ty7XEFT1wPrG1yB+YWOoRDQ1udTx8QUPPrbXW68UNJIvzifdDwd9rTu2a/j
PAuWULQGy3v02ynzapaJRYZUN6F+8RAiAQ1tPD61xK9GpNjs8ABh8/m0bBPuOXqr
+EaXb6dzxoo/mghH4PuKauAj7EIiTfi/uqRdIsz8pJatctFHqdaQrWw6CNR+AWCq
yxcCJbJZZBJJsSaDLu0lkmFx+NCENR8nKWW0FwL7jEGq3IdDAop4tia0dVAyFMS1
5H9aCMp1ThaMFpMvGrwgKYZyBDMePdy1/G+tM3HarPZVeVnsazFHBWe55VqjwcUH
9TsrL8L5Oxt234NA0aEVOzGrmL9cEmlqyAIxT18ixseZV9ucNiLEvrZaBZV3kx0n
J5ZiotUbtl7xc67IUweCPiT3TwlpPPExETkG1SGJJLRoYQrB1SaQ7LZkhEug29qx
77yAflGdsVa+6tF868gmy2yPvb8Xf5jugzXFPnxZDkMlbXgk137AwZesxuKIDAxE
G6ICFVWbDWxO73ou4jCDbry2ErqIAEXQRtPmzAMeXAf/7pwidwOXxQLY5N/+/FuY
Pt/I0Y0LaS83U0FkveFMSUgsBU8KGXK5GClIl448onATkz7ISA91pRholPH7DU4F
30qg/KlfDVBxNSAhMKWwDpdz/HEzCP5wn2Fe/Zr7tDzw/o/kgyc0CfONW8iK8AEj
vSyB3oNXPA8llAg4L80OrFS5jcI/p+QdoxIuqJlTtZjO23eZsXC95Uo+sgFHR8T+
JobZroncWFBp1Z3eTZN1utFoMB1mveDMINIvo2B/7WK5GAazyURwm++BpgMpfT/F
K1a/R3tXafr53kqGYqy3SoCJu428MrkF7Jiv74S5LtzNfw8LOSaWiXfrNOK72vR6
l4ZMPQXIUA9jNLVbUvywJuyne4jJ9tWBwXprqk1do31/4Nh1Cktr6FGHcS56W2Y/
qHzYH2pkM4bjfXA9UOy63obI52coyekyKQ7OTw6xmBuPhhvEET2ziRZVOwcSrLFq
ZzLr75xL/CPdz3Tsm1A06ZsWp6r8kiHLCFAbGI6XkA8sbdYaO23zPmD9OlQ+Zr3Q
TTw1H/H6QWWsn3vNJ/MMBTsjxyG2x/pVvNrALSD5cYnRDF6K+EFw1ld3g/LhiD9n
SC/RTglyxk1ZbqFvAH7NdE/vXrogW4w8N0ixkbYOKS0EqVpYiBj1DVcpkCJISDU4
RkxRFXMevffjqn5LqRK9+qcDiB4Oy2AygP6SO5K1qJGZzQa0wQRyEtICBTcMqKRp
dGa7PbFY3fXDOXGhnQcK2j0PheueSFQNpA/jipCI42pdP2vA88s2CJoNSTbKW3IR
jZBHyHNjjF/aWQzsAyC0QRM0AQe4H3Kq5I+ye2PXMR2uVUjM6ycCAeBZl/7lAIrt
6ERkDDgAsNxE6LHRxVR0BCPO7zuY/4On+UFMKyyRx+uyoEg6BmvrL0KkWx4REfv6
GNR5PzyDBE0MRnGV1ld6iFPaPdhtgXtMDF5DYgxTHV2uDiqogyQYGlBQ8rYiRmcy
fg53l3RFB2OH/vV+yc8BiM2tdY5a4EG8j31hmij5/N5tsb3Q3/97I8aRPIjMs/wV
qdcieZTI8IkHHGCtX/5dAp7BecYThUjg/cZBQ0UPFEjln3LF0JWxVZgO4s6YVNCa
dgyxmuqtMIsQA19IfnTNh8HXxZDtOSmjA5o/VWRuTxc1yfLzkFY+5hdqV80wSeke
fEfrgr3UczM/VZhCZr/HFNVjTRxLkZ5RJrxaV7a4AErEkeEFdTqgasc9OfbIuorW
hdk39L9H7ac9xiv9IqGJxgo+LHaFfbtpMMh0T6ZMVcC9o6y2k2Zt5W1A3iyb/e6+
5g6bkUoXpizvfiPDEOgCdoC3nFwFe761ORnmHbxpb7UCOuFulyhfRkIS/coD9pUD
jUY5JwcBqcz6wTFplwJcxwOzonhKz3h4qdOJqrIVJLRCcy7l9ALYQdSCW/4MKjy6
IUsT+x6tg14g15mJYhYFVcF9qjRd4zfI+J4Z81b5lTLiWK4Fs0Xgv28oIa5odFkV
mkTEZYm3ww1dHKwP2Lq7aF+ZkHYfZZOVlj1RBqBO8lkNYaV0NXsr31Kbk8gM/G9s
Yh6TFKTAnDLqxrjp2VrfCoGsPZzWg/6M8fjFlDMaecJEC88r7+GU3V2Rz103Da8w
yGMPKuGVFiDczwwyaSyIAa8WbjU2RdsqIjECD99S9srpgPLaZRQBzlquX8Toeycm
7OuneYdz9dYQy2HZM8kzxyl5JSK+hTvv2jye41H5McMQ8K0XlASNFFcM8R7Qf62v
TmTpJn1/zxH4xWD1Ne3CQWqeC7wwQVXqyNZCXc7SdtIxqVGi3BHXgTF7bhcgWtdZ
Eja5qiuNIPNu7RjmRK7WW0Lwf5F9zdQQPKP/UEGnZHb1SwbkzQlmkVadK9IC+Hsl
HV59FXcD1jYnxGMNINlf5Tq3itItQ95qbsFXjf0mN5o727N+hD9IqozcwcgUQlp1
P5ikCMdOE+JqCFO5q3XLJxilebxlS298G2Dz/C9AFjPkkhDZBiK8Qi43Ad6J+nV+
ZZ44yBugGTgOLsTBODXsLe5ERdoh+bGS2b5Th8CZofXW05k1t7eI7sqYy0iOUfUT
Vqs0nBPWic8VEt5Zk6/4H8fIhpriKEk1O/xr+vfp7eExoe/+MCQcVAUBaEcpZKLX
08ljpmXrZVd8OZkUTyyMaxFrKiULej1B4VOZWpbl5NWBCXZaRT4vEKqu0tvhsqs3
OuSHJJWYgqoCeegwpIKNr2Jcyal3oaw6rJ4QpanqGuOPc8JVamuPb2YD6l9jS12j
e0LTevJy34TdRJdjB2CwVl/L2d77s20Nm0c8B69RoFwk0+kNOkEimC8okZlSAzEo
331iLLaBYEu1VuvxxUMoBrAJ/ACUXWS/xji1k6trbJLx4ZkZWFCMuponx+phRGco
8CuBcnVaPikGOzLSTU2Efl4lfC2cPYWLVESiU64SOVlX2/CJPN66xbbr3SP24X6a
bCR6WY5Xaimvb3wgZ3owKZhQeHUEXOFqBgvjhp6KtFbwigVvas+4Zt4InZxFqYXO
wHiaEKVa7ppp9Zwxc4wM0gIjFtTPOdLAp2p8naQo5F8j+2Oe/Fj3LWXFLUl2fJOI
qOnnPqq/MlF8NbGOcMY1SLyEn4LdRM71gGvlrbdZMXKcFXPVjD5SRPtLgmzwivrX
2VDIwxiGcRzx1D2g/UOww16fB5ZlAVmBbxVeJI9RW9i3M8L5895wiieMKfKIkosg
TtXcLRq0JQ7hZc3w0sKCz1SLQoHACLNP1fKAfBNDyWm8jznmpnhaTDdOuOlqVaLi
ECAg99RTbdSBsu/6BM70n45KAs65x9a1LHaC9Cr2RiT+Nn0Giq6wpT4pUA5GWWm2
H5ZaVQao82ebQ8oWmiHQcGecFao5ZCXNCi8hjBStsFlsZI8ihafWep1+wJ5r4RqT
p6lGvoTtCS2fWjMgR403jBlLi2DzRB8jNeb8C9bBxDHzOMQ2yoxiRc4HUuOy9i4V
7w8KWQeeClT6B8DMJBo6tvXvimX9sIRjGhxpJbpGlNR3cdwvJcl7G0FG/ZpP+daz
Mie5Tekz4PvE4AXEVeDLcTwJ2C9HsmLxPTi4MmOhW6AmZo7ZC8LN2Ip4lPGBGCeV
NKfq3EbPBe6v4o7ejBe+mX+dgyX/cblpxUzklwu0M5/ErT0Mqvq+Rc2nI5xuExde
wNl+qoXNVFAjmqcCQJM0shYFvHtT/Mxl7OMDgeKHzRd2QtNHtP9D3lqsgm2eS585
fejIh7V0hPV4rFn+aGaHbWgpT6OKYRCoMOdXhBH7cJm3m23VTyr5EYZyJNeRWG/R
w9tQszWpzCWkobFxGanzcXvltA7gFP7rbzQTg94vjvNrBc/9rFaMCLtUMhuLE87J
fJRozJCrSCoAncdYZCUU2JquXGPJSpgegx5kBwuX/VFz4rItaE3EPFtlUHlqdh8s
yUVZN92NGHl/RPdRobwfjmaMlTFJkWu1kp7HnV2bO+89p1xuOOqoA/Wuv2j4IY0H
m+lj39U/4+8QBn4GR/VLrmauby45qeXzh1JMxLFjzWqEgCAU5SwHpjSpotEreV43
ECi3U+uOAwFWWuhjintWUaiSIc0SL4htsn2wgTqEmCLVL5x7sgxNf9jpGDSFD11z
QlsnsgeTj3O9vPYnfVO1vKc2jV3gWOQfLSZiEuMH0ATRXyDGbWh9U99mkoC1g9hE
0LQhY5G+NMblugEanuXF4GLo1WQyoxEL7VzZutdwFQRGjq5eg9CvFZkK0rVaXFNQ
MUNaO0+aTAtiahD7vKaCzoneoksS/EoQhNWvrzlrBi5ArYkWtPEY0p95la64kdjo
7QS7YKdhNiPV+9oPNBuGie3LKfaQRRfVc1sFIkdeQDc0jrXaLWaw9qjLwjpp/wip
AjeXN/ppteg4WUMWB65sxtiNJzDKwVCsRc4xAnImY3XAyecAuT8mzC4o/38oInmI
16Ilp5MMBNP9dDPUnWGC9SRwR1BIyk/biAUPFRktlFiCpDNA/EDZ870Mb/OaQz7w
GCtzkfiziv//YjR7v+5K+WA9wAO81e+MFusL1g5DxJywLYqwSoplLOtz+6E5lSQD
KTcN/dqzeOHxfp62/VIHz+wYu5m4tKrgoXYDO2IwMO1cdjR2MPml8LujkiQa7cgt
cY3SqSAhszAThSvj7/AGBhbDC/iSxjz6fYl6tLkr0JyPiv9anWKJcAK6QFzVdQj/
1YpglhGDKvn10idi5Cd0LWESzcplDRpYfVvS4qbHnjN219eL9QMzYweFfqN9FMdm
E4dv7hRVnoBK1SZaGHW0gta3+wLeK362dI4BjoyzZc7Bx5u5+2Vg6TUCHixDGYMI
AkCSML+aBAQ667KshkaVNCISsCE8x2fpUDqUASRFwokMeO9j2g74jJGIIsEZKhbf
kkkmJhioRWOAcAL4z7UuN+4LV5LNCRaljcRqL4/jfDN2bzWBamVl5Tw9pibKvsJn
wYvhyAq0EUGg5SWlnH6xyvljy1x+akwQUKyjGA+VyVXRnBVT/viBlzN5auF9Vvf8
sQIH6F9Afjhu8zwn22A1Y2icuuTNntA21gAZoAT4HJIreYN8xnTjBZVwKGM87nFr
/kfCv8DDMbymCvbuHqXi7T4rlghYP3QoYtYhFdXsfw2Das/Sq4Bt8E6u98YEMwI6
xdNGlwofwR1y8G5s7k+ZU1eksY3qNvZ4fts4H1STIWksNy5kksZFFVyQYKGX0A1m
4ZeyxX5SKV2EJ4K0XiIadBG4UY9ZJzE0RGs6iTK1AGGbXgv73ZyTsfWNp5u0kxCT
H4EYo92Ao30mVu62QqvJFnCqKsN7C0CGArdYabOKQba4gC3JgWo9dmwsdjKr17wt
lVWBQfNDFA5e0+FGujCqd6y4zHJgcZL44myjIhJdUEoIVgbI5mf/61E6hr6f/jJ4
pg0Fuit2u9c75t86ga+LUqBBLZ24OHXbo5VWKhN6dqrwEqBK+hWk10+9jG4pL3MB
Wtrtsm3a4m753ZsJE48n41vyiSB6nl7QvhggeCNFauynfRAqGlQVtnH9S6Oi4eRD
CkRu5KMup0270JZ3gZ/Pq8ljszgfuvf6g31qoyTYS4lAYDhW+WXdhnwHb1/hMClh
OriGw/JpJxFsLF4Bq98j+sG/2aPm5aCXEcuV1Sk2rrTvF5MFeNa2elJV5QfjRbj5
zeiv3Ayat9t9yMGEZfsI60xGPrfFIhaqGecI9rfQVkAoJPqO5gX5a8r/PE39o7yQ
boktUDMQ67pciAmMGu6bJCbw0JvTbtfJDfgMf9WRYo5o2RpgWul+zJVn2ePHGF5/
Sgko6jVz/RflH019GjSoDJIESsGPK/KPIY60PD6DcObF+FUAUwB+GNpIlyb6/KxR
gcfF2E3AadBTq/7sJ8UxrnAjSae3Koa0u2oMnpNh8iJrw1gVV+4ShyBzhguaERWA
Bm0kSBNHUoHSo7OMs9F8vfhWPdrn+r/djvfdLwJTQje6Xrmy1GzeLhG4ZSo1HGja
5QaWKJEh7nN/fx7yExZLLvJcdzkyiRsTImnbxs88RkNRyNT4MQEcN+yG0rRR1B6L
2FSmCOzykwVsf8eMlTvaWgM2dXcWrOOeUQjcZh64wLMpUTKL9oqpiLOzHTfXGZMi
YY7nfhHEeH0tmGZx9CYfDyo8/cfrGuJ1ufZePsRgGTKmjveaGL3gdDXlVXYfZdLu
uWIlLpZ5y9vKpjg/xUNsbirUnOPcyqnkiQaEyif5gS7GKxbtUhd4VPwAqPRFVUbd
DvTyNYJD6cp2oNi6eI+Iebv5sXX2IYu2+EsNo6rQ+oQMWbkprWhwYKaZ+LTnB0vm
YNuoJYi4WHWmnqaqe6mIdjl5dH3SGzdCfpjrbbRqZNhMDOs4JbJ8N9pGVSZzBBiV
DQOrTqGKrqTnJKo9SxKnx6IPgrRJnY50iL/YW9OW9e6UzJmn34Ipjp531Hb1/2TK
bfF5eWB5C0dkq8EJlVXGyZ8JgaQWupwf5fpuqi2zSRmd76ldND3tHuPBXzQq9YJ6
Z8hhiPqmhxGLLtzJ1pucMWvJFyD+6EzQ3i14cNyUdpe9HRr9Bbx3Ib+Bs8QSNfQS
zKxzYBpGZp6987re126OmIjx7+v+UiVys7HUfSFq3e/Rx6OqjY25sllAfCZTk7dT
jfkLFN2y1fkuDoFw3TEbUEEE6mq2jmbduPH/u3Yfd3PIT0mnzOOSp/34CeG0tdmt
U1atXJjrDkv8nlbI95EGvRJR5nrDbpfmMknTAfGYK32irZDyXQgeTC2gnL1mO8kq
83EeJ7gZ5q16WDeuGCXzLolghc92Mq8E6VqGcuAytt0HVxqJMgcxuJpHhl2bUtSa
EkQ9ZNbqPyLee0xjUPrnKwszuwUO2Hg2r3fcQyzcQIqtt0lv0SESF0aiFya/AMZ9
4PrkQLtOjMK7qt5+rYKetLLLGqNPFwirACCy4EUDUwuhu0MuBUBBh7vnnEzR6ZQn
xQ4lCHHL5j7Iai4AiM8qWaPMGgd0rn33DdXtzQv24maKYrsTK6TFytcYDyCS8KKF
cSRmLHSNiiIjHuXhBY3BWCTp8JEPGMzQgP9JEMWjPFWzwcc3gkTnN7rlERJ4slbv
wMqWiBe5j+IAd8ze9WB08/qC2Xun0k4DKiEzKd6m6rfqhYfqvdSXaUXlgnInki21
FyXCs2yKm6ojGZUOKp+4M2AChw6JRUPlytLPOe3eCh0j13ZrTx09Q12h+7nvZySY
iybot1yMrHp6PIx5LopeAnqFMNpUVAUzOFrROp2YGYcuDO9ajTwrtEzFki5uhnin
02MAn9TKNTVNRg/dn8myZtJJb4rC9E8PI1TKlu6LICRphrjOjtM1wm3pIRb0Kvk4
zIIrmxg9dj3a4vzkkC9m1PLbc6PYdDrweJQXEqBehYexoIiB86GZz9noCdIsvq1j
067RatDxM5iTvWve2hpLPS9AKfoTxFA7za61fDguCim/QOTXRaTbaS96Tl0K4JNt
474Yy8Dn4hym9wgKdYD1QSghi8Oy069lnc1TG/KlWJ8x46YCaTKE9vch98pt6qUo
Lv1sKln/ZudGCIm+f+90D3Lbjyxc9T26RFfnWLE18NgZccZMmIe8P9p++9I450Qc
VHU7Yyl6JJb/meBhbiOot0jX7qfUqAc54fixuYK3svKGtoOQt9pV+TmzqwtjVUHI
EOn+/XlpRUX/q4u4vcNnReoMAqxjx0vZZO2tG09tlNuIN9TuqKJorFR3LkzwetTU
MV4N7eeBp8TyjSun9UyU+Y/QZ5/KrlOt7fss2Rnaz1hBhCZoLcfDU6uObcOas7Sg
ZsI8s4RlrMaK25HWYeZ35dNwPLWlh7JrCnE1QscRcAxXvXdg0J2tzpFGBIc2TTWp
6XayvfoIJsnbBiKEjWmcSryLchZ6vcqDd49iqhpJ3XxTxLiET26z5Ryw4xU79zPq
NV6JrvWCGii6ikTc7IqMlEWertYFkmnoMcafvvNPwE+2ODx0nmk43xU7rNixz2/z
W4ls5tBUo0FV0XHHSNgBAqKJGIZ5WyfmmSoZ4VFUwnHqkKhCiy6f8QMSIh6L4gyD
fiP64uJbqxke7sPKdgqOwoBCgndW4H+gx/PHw3fiZDB3QgdVkqK7QU14lQTFDa1/
ibd9BsHLEXUZHhnR/4W/AZcG1oy1vHIr3sjKt3cRgFU26LjnAcCSLHpidyLI64iP
WwH8A5n97yXArfySf50ODcHQ3NFaeQGx2hk+SIpATeTtrBpRHuBppYILYNe7lXEa
J0u5y4B4yaieO937zCXXJE/pbLSrECh/Rrchu0B+SFrzfs7mgwaP775ZusK6pZ6A
X2XW5vKvcMDipxshGoAm2WRDIHi9GSKLB44VJZonuas4aZCHdJEvnbT7AeozsjLu
12ZvLLpc6vlIALWCtkTUw88kculKKj347kZSoaFpQSy4+KLQRwspD6jor/VkmZsY
sVg/RN6LCitJVygJ078hb/EPCy3z05Uydow+vt0k/w1TlG+7NeJcA8C+WubeGUZ/
snN9PW/Py1UO9o99jChP03flVuacDQHpRxdIX98j1HJucrNttjGs1GCBeDqfaFap
jJIqK/gz4CH6AqhgZHvvnJuPdupKouQmwhiX3UpC4DX09ueqQo/C6IGYDeRZfo9b
/xe8DOmi601adap1y31zT7dv7SpQrz2DbWjLY/ZLdDxJKGA2GnZHsjyEs5L7epsz
bHXtbIHauztpMKypQgSdqD57zEf2o6ySk0qO3uyKFYd22XzqEAtkJ510uPDzjyIo
/9GMpj3tRPffN9c7K1cGK6iMPDcs7RtE7wDmB2aSeHjkehQl4DF5MM3RQJMmhD6J
JHkA59uaTbKT6zOOi6hr0tEAS84DrwjRpc/UQ9GG/y7ZcRgPeOVWf8sKVAbEs4Bp
Uw9l0NQtL+Hzs9PW4oAgaLTc4nWs8IaZdOxMRzRM2Fn7O6B9Xx7b2VwrhBu5tmku
GdRATClnIrSgaeZr/xTdvTuEA3j8M6ApudExzHOrpx08z91ZJ590ObtOe+kc+YRk
vtB+QfuK3CZmTqK5BY+qNRuVLWzVp80VXFejFIUacVnY2j3/pFM3t1Tijv/QYvyn
56hhDsPtAELALKxaT914MjHskBlNKzJmqZAPV8wIm20EIeJZzaaTbtN9g10LVj/O
JksiSNDtLimHru2GOgG54YSdIOPjr0CLLLmnyiX88i6uezscEix5OETQJq88GYA0
W/CQJnMeNNZzTjHQhKHU2dIHO6hM0cB8e+mVYea06xO57x/7ErIGFs6Vh/DAz5w/
1ZXGSnxpK40dClQdjUPJyBHGlYs4vPxz1HUaZnFn6jAT/Ai4ZxoQL8aVmlVWW9PM
vb6Cj3wH9db6GIsakawxLLp274xxWyg4llKCZD1joW9481570iIKkysweB6Qzbe8
3RQfaeIPX0xsgPLqGjSIfyZEoCwpMe4Hz2lRThvsDKiUnVq+Pq5vO4F2NhP/Hjdv
30oQ7Yvx1YXzYD1fUo113MiQHIkF7K9z3F3FYqyi8ZvGxlhaoksSE41sEOVqVeXd
O9GgIg5xclC5Yp62085jeeDrZRZmZwd7rnqjPIH+S22oy+O6/WZ+FvFH0n5CDQ93
g4glz4QBqi8OPJaUjr7ooAWDUqJrpGQO62weaQJlmcgbbSR78EZ4p3Dv4rt6WGGv
lCEFFWNQxaUSGuco/GGjTNzUsBoQ3ZmZbh0JBLbw7Rtx3tgUH7WtTijZG7aaOxG2
TXH7XBQsFmn7LmAI2pAnPheW8noe3x/gRtDkAczJmE2cMcli4supQ2yRtHx/vnpK
qdmGg6yONk0uq9yhsmbiMf/g73qTa+pp9UpF1QEIeOADPO1DgSmQVDpz/Guxe+MR
+kdihkzjMuSm37SyesbCBe8cYEj00RhlY2Op8Ye4cBbAhzk0jwwCea2KXpjdiCBg
u9pcnNiDm1GRPTqeHsS6bFyfPsb7avJZ3Bb9GdxQ+T85rRm6CJIoHlhbiC+C4tUu
RtHh6r6m8D9tOlziLjvn/cCykWGHcArXImFlPuhHztfan/hkud+mr8BgGcVX6pR6
ZFs/gi04AUfsNyS+sfCrLV2zbB7xzJ+1okWyBMbxyEzwXbe+7z3iO2wvjmaRqOZa
j+Hpv820nTBItZ+AsXfTbA4h6xCKYUr7jZNvBOdNph7jF8Ic/Ok4pQ6xSkpZHJDF
wM/JPcFapcSn/2hnOYVsORmgBIQ3iTzwFhSIGJxN1h1OWC5DXmNsEEeHBt3HLCOI
j9IZcPndvrM5zp1/jnAMUEHVTLmq9CWnQ/RPKpYVCZoQ/nB+OMMRz6ap2+MJtva0
zQmixHDBrn+fooZzqmv34vpoqP0LHoxQqUn/wJaG6s9ZP8oAeD9OPbX8vI4wvvwS
tTvEo6Zsgtu0+T4KrEKn6+HxtI53hhgCiJxYwL+DrfBCwVR00jFbRkVDqBHDskIJ
MFUoFK+p0EDm/gTe+Qp0/iNh/OQhN8FNG8ETtTv849oe5xK1gtaaACpA/wV1if2w
Qy8m7CfJ/gxKURRxXz5+juHVskpRGnUUFLDVANM6QhSmcxu3pNP625csbttC06Ah
CLhNknni2psOH9wlbICjmLjz+8apVuQoVyrmPSvmNOoOlsPs81bz349JKSQXTnil
4M9+rWnU0u0oXq66ykL1UDZSD0B/MNdAnMDVzzG1BFudUOkwehnkxd4edQzXRkES
yOpUzBiLZIebEY5B9i+M0MKvyWtwLhVuOcH+Uj4gpql6gmGLM4fiXu0JRSaQqJ9b
X3eXCte+tVXAL1uLgU+zRD6qrfjxT4eHDApscPFWdHi+o1z5Q6lSMtAPugPXoQR9
qxxB0XsRTtyRC2CAYP/xiVdr24qNwD5it/qsvGO+RgNY1fZ0hzC/iEizv17deCzs
8+6EPB/G6e1aoUAWCndYsGltaeBc2rIHgTy8S+JVZP9wghLCaEZE94SuxeEcBsFK
+tqGP/h6woQ5kw1AwgkT66UExEQe+Volv1WdCurtLZRGL/hNxG65qw+0nGfRGs4f
q952wG76CvDMegCj0q+iceXjwGNYuclmq3R5S2xOq9kVd9WdEL1FoeWLilWxu0mC
yBAmYD9kG9OMhKZQsjJGJuo3ZU/VLddPcGtGKQU2ZV3QASpm94II2Vb21RqqIS6i
H3Qqfuo2+Y+2gsppfzCrpiGRnGQRJQtDpb7x4LUfvZx/TkaH2k01dzyP6freva5F
758gcbMFImNZkCrtXwhKaKu0mHcrVqWdJXuxkFO9TqpydOb9oLbsRmOg9XbAWkVa
GV4Ju4VJxGX0kOPdPgdo6MXtVdsPwy34j+IZTbSlekZvGt/WNC8vBEnofoC/9whG
2rFIZQQvEeTYbDoYDveea7geJfh3w1CUm3+CCn24vrlmWEEEjFvFD7BaF3sEPBj+
veSJGOLrNrmU0Bml2B2sxdj1B8mACV4fr8vlTlM+BCcfeVC3nMdrzwrRAJtMGpWS
cZDr1TRpcQTsaWyrIzCvhXb4wCVhqWfjkghhNLiEEO1jp70SCk0E7UYxcTev0gvR
/7XLkbFUt77k5Ms3M1Hkr50GIZnGIdnGfEyV+osdRPS/D3/r2P63YvnNKPA6SFSU
K8MKRTNlm2kbYRVmEiJmMvY7WyfIsmRBEG5aeEfOg8RLssT/L8l/nBlJyFeFfV91
PMxEUmsxwqs374AK8Mt9y8nSter63tjUu5ffNZadf5AyDdqj2mggWLdS3ZVwwabp
09xn+1YdfbKeCsY16Amn0P57lX2695suqLB8Y/Zmf1fsyJlaOwJ7YlaoAsTt9Xrw
6o3QEwXuiuZeN+xE4Bc2jA2aaMVvnUJrFgxE6lPzTSQ4r85jFnZN8yu7H4RtZyQd
nRJd0OrDNgolzpd7LiWDryEJt9OSJ7U3R2RAcOO9GFb3ID8T88BewJhbe0xpU4Cs
Bg1Ou6IMDWC6CiFtv0PJFbnm+RCr5ftls8bgtX6DN7NfDHkmDFiD3rphx2612jmc
t8+lONITTe3g+RSIISsLgeApVIBPKejD7ZDPLtE0CWuQZ5sVwgWlR3bNUaytqw7+
`pragma protect end_protected

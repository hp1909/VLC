module delay(
	input	[31:0] iData,
	output	[31:0] oData
	);
assign oData =iData;
endmodule